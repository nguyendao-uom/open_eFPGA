##
## LEF for PtnCells ;
## created by Innovus v19.11-s128_1 on Mon Dec  6 14:59:22 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO E_CPU_IO_bot
  CLASS BLOCK ;
  SIZE 200.100000 BY 200.260000 ;
  FOREIGN E_CPU_IO_bot 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3908 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.846 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.80613 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.6559 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 9.240000 0.000000 9.620000 0.700000 ;
    END
  END N1END[3]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.859 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.56801 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 10.4653 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 7.860000 0.000000 8.240000 0.700000 ;
    END
  END N1END[2]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3194 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.489 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.74606 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.9529 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 6.480000 0.000000 6.860000 0.700000 ;
    END
  END N1END[1]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.353 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.657 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.94141 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.3259 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 0.000000 5.480000 0.700000 ;
    END
  END N1END[0]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.933 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.439 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.91111 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 28.0155 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 21.660000 0.000000 22.040000 0.700000 ;
    END
  END N2MID[7]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4786 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.285 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 15.0543 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 73.8902 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 19.820000 0.000000 20.200000 0.700000 ;
    END
  END N2MID[6]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.033 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.057 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 15.4389 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 75.8135 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 18.440000 0.000000 18.820000 0.700000 ;
    END
  END N2MID[5]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9818 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.683 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.91946 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.05724 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 17.060000 0.000000 17.440000 0.700000 ;
    END
  END N2MID[4]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3834 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.809 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 14.9858 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 72.1515 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 15.680000 0.000000 16.060000 0.700000 ;
    END
  END N2MID[3]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9858 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.821 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 14.8242 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 72.7401 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 13.840000 0.000000 14.220000 0.700000 ;
    END
  END N2MID[2]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9164 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.464 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.22094 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.7165 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 12.460000 0.000000 12.840000 0.700000 ;
    END
  END N2MID[1]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1445 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.0218 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.92 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 27.1392 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 142.409 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 11.080000 0.000000 11.460000 0.700000 ;
    END
  END N2MID[0]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.027 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.85933 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 16.763 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 33.620000 0.000000 34.000000 0.700000 ;
    END
  END N2END[7]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.88 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.58673 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.5589 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 32.240000 0.000000 32.620000 0.700000 ;
    END
  END N2END[6]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.605 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.917 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.91246 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 48.1811 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 30.860000 0.000000 31.240000 0.700000 ;
    END
  END N2END[5]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3194 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.489 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.8499 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.8747 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 29.020000 0.000000 29.400000 0.700000 ;
    END
  END N2END[4]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2234 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.009 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 16.1712 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 78.3764 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 27.640000 0.000000 28.020000 0.700000 ;
    END
  END N2END[3]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9985 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.8315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.1938 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 26.2318 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 138.494 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 26.260000 0.000000 26.640000 0.700000 ;
    END
  END N2END[2]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6998 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.391 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 15.2485 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 74.8613 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 24.420000 0.000000 24.800000 0.700000 ;
    END
  END N2END[1]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6569 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.2048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.896 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 26.497 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 140.458 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 23.040000 0.000000 23.420000 0.700000 ;
    END
  END N2END[0]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.441 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.979 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.62465 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 11.5832 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 58.000000 0.000000 58.380000 0.700000 ;
    END
  END N4END[15]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.1318 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.84 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 10.9609 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 56.2761 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 56.620000 0.000000 57.000000 0.700000 ;
    END
  END N4END[14]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.837 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.82397 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.67071 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 54.780000 0.000000 55.160000 0.700000 ;
    END
  END N4END[13]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.755 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.2202 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.402 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 53.400000 0.000000 53.780000 0.700000 ;
    END
  END N4END[12]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1849 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.1908 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.488 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 25.9487 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 137.077 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 52.020000 0.000000 52.400000 0.700000 ;
    END
  END N4END[11]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5858 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.703 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.28956 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.9987 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 50.180000 0.000000 50.560000 0.700000 ;
    END
  END N4END[10]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7208 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.496 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 11.8263 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 57.7502 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 48.800000 0.000000 49.180000 0.700000 ;
    END
  END N4END[9]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.1568 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.64 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 12.2137 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 61.7549 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 47.420000 0.000000 47.800000 0.700000 ;
    END
  END N4END[8]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.871 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 14.5548 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 70.1017 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 45.580000 0.000000 45.960000 0.700000 ;
    END
  END N4END[7]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5826 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.687 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.63205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.7111 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 44.200000 0.000000 44.580000 0.700000 ;
    END
  END N4END[6]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 11.8483 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 56.464 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 42.820000 0.000000 43.200000 0.700000 ;
    END
  END N4END[5]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7952 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.75 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.16801 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.604 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 41.440000 0.000000 41.820000 0.700000 ;
    END
  END N4END[4]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5357 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.5175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.5448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.376 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 36.2171 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 191.363 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 39.600000 0.000000 39.980000 0.700000 ;
    END
  END N4END[3]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7175 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.1148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 30.5183 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 159.644 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 38.220000 0.000000 38.600000 0.700000 ;
    END
  END N4END[2]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.837 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.01872 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.5535 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 36.840000 0.000000 37.220000 0.700000 ;
    END
  END N4END[1]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1521 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.3248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 135.536 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 37.3952 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 197.512 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 35.000000 0.000000 35.380000 0.700000 ;
    END
  END N4END[0]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8698 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.123 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.87354 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 12.8276 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 82.380000 0.000000 82.760000 0.700000 ;
    END
  END NN4END[15]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6944 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.311 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.2928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.032 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 12.4051 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 62.6714 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 80.540000 0.000000 80.920000 0.700000 ;
    END
  END NN4END[14]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.775 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.96215 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.3616 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 79.160000 0.000000 79.540000 0.700000 ;
    END
  END NN4END[13]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5906 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 10.842 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 52.829 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 77.780000 0.000000 78.160000 0.700000 ;
    END
  END NN4END[12]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2733 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.9106 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.464 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 21.2591 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 111.797 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 75.940000 0.000000 76.320000 0.700000 ;
    END
  END NN4END[11]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3649 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9498 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.536 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 18.3345 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 96.7448 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 74.560000 0.000000 74.940000 0.700000 ;
    END
  END NN4END[10]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.9708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.648 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 10.7488 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 55.6646 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 73.180000 0.000000 73.560000 0.700000 ;
    END
  END NN4END[9]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9565 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.1796 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 119.232 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 32.7274 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 173.395 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 71.800000 0.000000 72.180000 0.700000 ;
    END
  END NN4END[8]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8906 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.345 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 13.4521 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 65.8296 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 69.960000 0.000000 70.340000 0.700000 ;
    END
  END NN4END[7]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5963 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.8468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.32 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 17.1026 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 88.2034 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 68.580000 0.000000 68.960000 0.700000 ;
    END
  END NN4END[6]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.837 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.82397 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.67071 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 67.200000 0.000000 67.580000 0.700000 ;
    END
  END NN4END[5]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.3716 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.256 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 27.6333 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 146.664 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 65.360000 0.000000 65.740000 0.700000 ;
    END
  END NN4END[4]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.5285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.1448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 21.1731 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 108.284 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 63.980000 0.000000 64.360000 0.700000 ;
    END
  END NN4END[3]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1693 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.7638 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 148.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 39.9352 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 211.308 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 62.600000 0.000000 62.980000 0.700000 ;
    END
  END NN4END[2]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2795 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.2365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.7818 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 116.64 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 31.0773 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 164.333 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 60.760000 0.000000 61.140000 0.700000 ;
    END
  END NN4END[1]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.774 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.19205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 9.56566 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 59.380000 0.000000 59.760000 0.700000 ;
    END
  END NN4END[0]
  PIN Ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.260000 0.000000 164.640000 0.700000 ;
    END
  END Ci
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 3.39138 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 15.6956 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 80.720000 0.700000 81.100000 ;
    END
  END E1END[3]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.392 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 2.89818 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 13.8586 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 79.500000 0.700000 79.880000 ;
    END
  END E1END[2]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 1.93764 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 8.22222 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 77.670000 0.700000 78.050000 ;
    END
  END E1END[1]
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.488 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 5.25468 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 26.2801 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 76.450000 0.700000 76.830000 ;
    END
  END E1END[0]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 92.920000 0.700000 93.300000 ;
    END
  END E2MID[7]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 3.33239 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 16.0202 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 91.090000 0.700000 91.470000 ;
    END
  END E2MID[6]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 2.36 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 10.334 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 89.870000 0.700000 90.250000 ;
    END
  END E2MID[5]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 88.040000 0.700000 88.420000 ;
    END
  END E2MID[4]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 86.820000 0.700000 87.200000 ;
    END
  END E2MID[3]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 3.08162 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 14.8498 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 84.990000 0.700000 85.370000 ;
    END
  END E2MID[2]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 1.97535 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 8.41077 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 83.770000 0.700000 84.150000 ;
    END
  END E2MID[1]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 81.940000 0.700000 82.320000 ;
    END
  END E2MID[0]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 104.510000 0.700000 104.890000 ;
    END
  END E2END[7]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 2.32983 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 10.3879 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 103.290000 0.700000 103.670000 ;
    END
  END E2END[6]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 2.02923 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 8.85926 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 101.460000 0.700000 101.840000 ;
    END
  END E2END[5]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 100.240000 0.700000 100.620000 ;
    END
  END E2END[4]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 98.410000 0.700000 98.790000 ;
    END
  END E2END[3]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 2.51293 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 10.0121 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 97.190000 0.700000 97.570000 ;
    END
  END E2END[2]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 2.32148 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 10.4081 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 95.360000 0.700000 95.740000 ;
    END
  END E2END[1]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 94.140000 0.700000 94.520000 ;
    END
  END E2END[0]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 128.300000 0.700000 128.680000 ;
    END
  END EE4END[15]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 127.080000 0.700000 127.460000 ;
    END
  END EE4END[14]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 125.250000 0.700000 125.630000 ;
    END
  END EE4END[13]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 124.030000 0.700000 124.410000 ;
    END
  END EE4END[12]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 122.200000 0.700000 122.580000 ;
    END
  END EE4END[11]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 120.980000 0.700000 121.360000 ;
    END
  END EE4END[10]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 119.150000 0.700000 119.530000 ;
    END
  END EE4END[9]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 117.930000 0.700000 118.310000 ;
    END
  END EE4END[8]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 116.710000 0.700000 117.090000 ;
    END
  END EE4END[7]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 114.880000 0.700000 115.260000 ;
    END
  END EE4END[6]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 113.660000 0.700000 114.040000 ;
    END
  END EE4END[5]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 111.830000 0.700000 112.210000 ;
    END
  END EE4END[4]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 110.610000 0.700000 110.990000 ;
    END
  END EE4END[3]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 108.780000 0.700000 109.160000 ;
    END
  END EE4END[2]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 107.560000 0.700000 107.940000 ;
    END
  END EE4END[1]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 105.730000 0.700000 106.110000 ;
    END
  END EE4END[0]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 73.8194 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 357.857 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.477381 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 145.990000 0.700000 146.370000 ;
    END
  END E6END[11]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 28.0619 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 127.601 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 144.770000 0.700000 145.150000 ;
    END
  END E6END[10]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 20.3417 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 89.5496 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 143.550000 0.700000 143.930000 ;
    END
  END E6END[9]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 17.4492 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 73.7044 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 141.720000 0.700000 142.100000 ;
    END
  END E6END[8]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 15.119 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 61.6329 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 140.500000 0.700000 140.880000 ;
    END
  END E6END[7]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9828 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 29.4143 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 141.097 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 138.670000 0.700000 139.050000 ;
    END
  END E6END[6]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.9146 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 191.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 29.1964 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 146.06 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 137.450000 0.700000 137.830000 ;
    END
  END E6END[5]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.8116 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 148.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 29.6004 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.508 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.636111 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 135.620000 0.700000 136.000000 ;
    END
  END E6END[4]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4752 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 33.3718 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 166.05 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 134.400000 0.700000 134.780000 ;
    END
  END E6END[3]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 21.9813 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 98.2163 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 132.570000 0.700000 132.950000 ;
    END
  END E6END[2]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.9146 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 191.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 21.1548 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 100.712 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 131.350000 0.700000 131.730000 ;
    END
  END E6END[1]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 88.4893 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 431.389 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.477381 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 130.130000 0.700000 130.510000 ;
    END
  END E6END[0]
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3458 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.503 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 88.360000 0.000000 88.740000 0.700000 ;
    END
  END S1BEG[3]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0185 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.3068 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.44 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 86.520000 0.000000 86.900000 0.700000 ;
    END
  END S1BEG[2]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.595 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.749 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 85.140000 0.000000 85.520000 0.700000 ;
    END
  END S1BEG[1]
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4861 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.0108 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.528 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 83.760000 0.000000 84.140000 0.700000 ;
    END
  END S1BEG[0]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.741 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 112.740000 0.000000 113.120000 0.700000 ;
    END
  END S2BEG[7]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7742 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.645 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 110.900000 0.000000 111.280000 0.700000 ;
    END
  END S2BEG[6]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9858 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.821 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 109.520000 0.000000 109.900000 0.700000 ;
    END
  END S2BEG[5]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3666 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 108.140000 0.000000 108.520000 0.700000 ;
    END
  END S2BEG[4]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.837 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 106.300000 0.000000 106.680000 0.700000 ;
    END
  END S2BEG[3]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0806 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.295 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 104.920000 0.000000 105.300000 0.700000 ;
    END
  END S2BEG[2]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5358 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.453 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 103.540000 0.000000 103.920000 0.700000 ;
    END
  END S2BEG[1]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3858 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.821 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 101.700000 0.000000 102.080000 0.700000 ;
    END
  END S2BEG[0]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.9828 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.712 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 100.320000 0.000000 100.700000 0.700000 ;
    END
  END S2BEGb[7]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7642 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.713 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 98.940000 0.000000 99.320000 0.700000 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7857 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.1888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.144 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 97.560000 0.000000 97.940000 0.700000 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3786 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.667 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 95.720000 0.000000 96.100000 0.700000 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3194 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.489 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 94.340000 0.000000 94.720000 0.700000 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6526 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.155 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 92.960000 0.000000 93.340000 0.700000 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2982 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.265 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 91.120000 0.000000 91.500000 0.700000 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9646 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.597 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 89.740000 0.000000 90.120000 0.700000 ;
    END
  END S2BEGb[0]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.335 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 136.660000 0.000000 137.040000 0.700000 ;
    END
  END S4BEG[15]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9174 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.361 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 135.280000 0.000000 135.660000 0.700000 ;
    END
  END S4BEG[14]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.527 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 133.900000 0.000000 134.280000 0.700000 ;
    END
  END S4BEG[13]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5574 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.679 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 132.060000 0.000000 132.440000 0.700000 ;
    END
  END S4BEG[12]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.441 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 130.680000 0.000000 131.060000 0.700000 ;
    END
  END S4BEG[11]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.955 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.667 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 129.300000 0.000000 129.680000 0.700000 ;
    END
  END S4BEG[10]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6522 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.153 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 127.460000 0.000000 127.840000 0.700000 ;
    END
  END S4BEG[9]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.907 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 126.080000 0.000000 126.460000 0.700000 ;
    END
  END S4BEG[8]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.599 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 124.700000 0.000000 125.080000 0.700000 ;
    END
  END S4BEG[7]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9238 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.511 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 123.320000 0.000000 123.700000 0.700000 ;
    END
  END S4BEG[6]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.419 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 121.480000 0.000000 121.860000 0.700000 ;
    END
  END S4BEG[5]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.129 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.537 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 120.100000 0.000000 120.480000 0.700000 ;
    END
  END S4BEG[4]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.9488 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.864 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 118.720000 0.000000 119.100000 0.700000 ;
    END
  END S4BEG[3]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.871 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 116.880000 0.000000 117.260000 0.700000 ;
    END
  END S4BEG[2]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.251 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 115.500000 0.000000 115.880000 0.700000 ;
    END
  END S4BEG[1]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.741 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 114.120000 0.000000 114.500000 0.700000 ;
    END
  END S4BEG[0]
  PIN SS4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.871 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 161.040000 0.000000 161.420000 0.700000 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3666 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 159.660000 0.000000 160.040000 0.700000 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1766 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.775 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.820000 0.000000 158.200000 0.700000 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.893 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.357 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 156.440000 0.000000 156.820000 0.700000 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5574 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.679 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 155.060000 0.000000 155.440000 0.700000 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.912 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.452 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 153.680000 0.000000 154.060000 0.700000 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4618 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.201 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 151.840000 0.000000 152.220000 0.700000 ;
    END
  END SS4BEG[9]
  PIN SS4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.067 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.227 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.460000 0.000000 150.840000 0.700000 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.241 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.097 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 149.080000 0.000000 149.460000 0.700000 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.585 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 147.240000 0.000000 147.620000 0.700000 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.784 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 145.860000 0.000000 146.240000 0.700000 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1766 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.775 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 144.480000 0.000000 144.860000 0.700000 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4882 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.215 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 142.640000 0.000000 143.020000 0.700000 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.741 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 141.260000 0.000000 141.640000 0.700000 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3222 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.503 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 139.880000 0.000000 140.260000 0.700000 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.907 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 138.500000 0.000000 138.880000 0.700000 ;
    END
  END SS4BEG[0]
  PIN W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.9654 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.144 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 9.350000 0.700000 9.730000 ;
    END
  END W1BEG[3]
  PIN W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 7.520000 0.700000 7.900000 ;
    END
  END W1BEG[2]
  PIN W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.2074 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 6.300000 0.700000 6.680000 ;
    END
  END W1BEG[1]
  PIN W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9513 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.872 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.4998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.136 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 5.080000 0.700000 5.460000 ;
    END
  END W1BEG[0]
  PIN W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.1144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.272 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 20.940000 0.700000 21.320000 ;
    END
  END W2BEG[7]
  PIN W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6836 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.2838 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 97.984 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 19.720000 0.700000 20.100000 ;
    END
  END W2BEG[6]
  PIN W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 17.890000 0.700000 18.270000 ;
    END
  END W2BEG[5]
  PIN W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.4944 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.632 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 16.670000 0.700000 17.050000 ;
    END
  END W2BEG[4]
  PIN W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.5304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.824 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 15.450000 0.700000 15.830000 ;
    END
  END W2BEG[3]
  PIN W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.2748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.336 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 13.620000 0.700000 14.000000 ;
    END
  END W2BEG[2]
  PIN W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 12.400000 0.700000 12.780000 ;
    END
  END W2BEG[1]
  PIN W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.6894 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.672 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 10.570000 0.700000 10.950000 ;
    END
  END W2BEG[0]
  PIN W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.712 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 33.140000 0.700000 33.520000 ;
    END
  END W2BEGb[7]
  PIN W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3046 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.5038 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 93.824 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 31.310000 0.700000 31.690000 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 30.090000 0.700000 30.470000 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 28.870000 0.700000 29.250000 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.1074 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.568 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 27.040000 0.700000 27.420000 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9256 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.4448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 120.176 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 25.820000 0.700000 26.200000 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 23.990000 0.700000 24.370000 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.5414 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.216 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 22.770000 0.700000 23.150000 ;
    END
  END W2BEGb[0]
  PIN WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 56.930000 0.700000 57.310000 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 55.100000 0.700000 55.480000 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 53.880000 0.700000 54.260000 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 52.660000 0.700000 53.040000 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 50.830000 0.700000 51.210000 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 49.610000 0.700000 49.990000 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 47.780000 0.700000 48.160000 ;
    END
  END WW4BEG[9]
  PIN WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.3684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.96 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 46.560000 0.700000 46.940000 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 44.730000 0.700000 45.110000 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 43.510000 0.700000 43.890000 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 42.290000 0.700000 42.670000 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 40.460000 0.700000 40.840000 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 39.240000 0.700000 39.620000 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 37.410000 0.700000 37.790000 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.2644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.072 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 36.190000 0.700000 36.570000 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 34.360000 0.700000 34.740000 ;
    END
  END WW4BEG[0]
  PIN W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.2644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.072 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 74.620000 0.700000 75.000000 ;
    END
  END W6BEG[11]
  PIN W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 73.400000 0.700000 73.780000 ;
    END
  END W6BEG[10]
  PIN W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.3004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.264 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 71.570000 0.700000 71.950000 ;
    END
  END W6BEG[9]
  PIN W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 70.350000 0.700000 70.730000 ;
    END
  END W6BEG[8]
  PIN W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.5064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.696 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 68.520000 0.700000 68.900000 ;
    END
  END W6BEG[7]
  PIN W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 67.300000 0.700000 67.680000 ;
    END
  END W6BEG[6]
  PIN W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 66.080000 0.700000 66.460000 ;
    END
  END W6BEG[5]
  PIN W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 64.250000 0.700000 64.630000 ;
    END
  END W6BEG[4]
  PIN W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.4744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.192 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 63.030000 0.700000 63.410000 ;
    END
  END W6BEG[3]
  PIN W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.3004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.264 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 61.200000 0.700000 61.580000 ;
    END
  END W6BEG[2]
  PIN W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 59.980000 0.700000 60.360000 ;
    END
  END W6BEG[1]
  PIN W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.3004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.264 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 58.150000 0.700000 58.530000 ;
    END
  END W6BEG[0]
  PIN OPA_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7796 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 17.356 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 85.1647 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 91.700000 200.100000 92.080000 ;
    END
  END OPA_I0
  PIN OPA_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 29.1246 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 139.712 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 94.750000 200.100000 95.130000 ;
    END
  END OPA_I1
  PIN OPA_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.5386 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 114.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 12.9742 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 61.4306 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 97.800000 200.100000 98.180000 ;
    END
  END OPA_I2
  PIN OPA_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 11.8571 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 46.6885 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.566667 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 100.240000 200.100000 100.620000 ;
    END
  END OPA_I3
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.002 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.608 LAYER met2  ;
    ANTENNAMAXAREACAR 1.13673 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 4.92502 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0299696 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 162.420000 0.000000 162.800000 0.700000 ;
    END
  END UserCLK
  PIN OPB_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 80.7905 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 391.288 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 80.110000 200.100000 80.490000 ;
    END
  END OPB_I0
  PIN OPB_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.52 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 17.2337 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 77.0933 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 83.160000 200.100000 83.540000 ;
    END
  END OPB_I1
  PIN OPB_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 24.3524 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 108.407 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 85.600000 200.100000 85.980000 ;
    END
  END OPB_I2
  PIN OPB_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.5866 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 115.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 17.7036 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 84.1806 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 88.650000 200.100000 89.030000 ;
    END
  END OPB_I3
  PIN RES0_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 68.520000 200.100000 68.900000 ;
    END
  END RES0_O0
  PIN RES0_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 71.570000 200.100000 71.950000 ;
    END
  END RES0_O1
  PIN RES0_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 74.010000 200.100000 74.390000 ;
    END
  END RES0_O2
  PIN RES0_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 77.060000 200.100000 77.440000 ;
    END
  END RES0_O3
  PIN RES1_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 56.930000 200.100000 57.310000 ;
    END
  END RES1_O0
  PIN RES1_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.5374 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.528 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 59.370000 200.100000 59.750000 ;
    END
  END RES1_O1
  PIN RES1_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 62.420000 200.100000 62.800000 ;
    END
  END RES1_O2
  PIN RES1_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 65.470000 200.100000 65.850000 ;
    END
  END RES1_O3
  PIN RES2_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 45.340000 200.100000 45.720000 ;
    END
  END RES2_O0
  PIN RES2_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 47.780000 200.100000 48.160000 ;
    END
  END RES2_O1
  PIN RES2_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 50.830000 200.100000 51.210000 ;
    END
  END RES2_O2
  PIN RES2_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 53.880000 200.100000 54.260000 ;
    END
  END RES2_O3
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 4.5209 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 199.560000 5.480000 200.260000 ;
    END
  END UserCLKo
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 37.5894 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 200.472 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 55.8124 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 290.417 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 194.180000 0.700000 194.560000 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 38.8158 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 192.377 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 192.350000 0.700000 192.730000 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 40.9464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 218.376 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 57.7747 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 302.583 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 191.130000 0.700000 191.510000 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 16.0476 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 78.6807 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 189.300000 0.700000 189.680000 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.6004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.864 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 27.1937 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 138.576 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 188.080000 0.700000 188.460000 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 14.8241 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 72.7659 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 186.250000 0.700000 186.630000 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 15.5171 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 73.8672 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 185.030000 0.700000 185.410000 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.96 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 17.8683 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 89.0152 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 183.200000 0.700000 183.580000 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 15.721 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 76.9288 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 181.980000 0.700000 182.360000 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.9344 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 170.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 53.2991 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 275.603 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 180.760000 0.700000 181.140000 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 15.4985 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 73.774 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 178.930000 0.700000 179.310000 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 12.3242 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 60.139 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 177.710000 0.700000 178.090000 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.9895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 192.88 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 76.0771 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 390.209 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 175.880000 0.700000 176.260000 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.92 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 23.852 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 115.8 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 174.660000 0.700000 175.040000 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.2004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.064 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 90.6028 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 452.812 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.50915 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 172.830000 0.700000 173.210000 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.0344 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 277.512 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 73.3054 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 381.875 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 171.610000 0.700000 171.990000 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 62.0345 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 305.756 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.50915 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 169.780000 0.700000 170.160000 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 19.6127 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 94.2032 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 168.560000 0.700000 168.940000 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.512 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 63.8522 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 317.426 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.50915 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 167.340000 0.700000 167.720000 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 51.2115 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 252.17 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 165.510000 0.700000 165.890000 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 7.15293 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 33.6795 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 164.290000 0.700000 164.670000 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 15.0418 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 73.7886 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 162.460000 0.700000 162.840000 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.92 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 5.9437 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 28.8458 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 161.240000 0.700000 161.620000 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 43.1748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 230.736 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 63.6058 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 336.579 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 159.410000 0.700000 159.790000 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.4584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 242.44 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 66.7028 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 352.54 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 158.190000 0.700000 158.570000 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 5.89185 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 27.8842 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 156.360000 0.700000 156.740000 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 19.9842 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 98.2842 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 155.140000 0.700000 155.520000 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 30.7548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 164.496 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 47.1467 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 248.64 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 153.920000 0.700000 154.300000 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 9.46377 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 44.7461 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 152.090000 0.700000 152.470000 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.736 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 15.223 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 76.9872 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 150.870000 0.700000 151.250000 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 15.1357 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 73.0599 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 149.040000 0.700000 149.420000 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.96 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 35.4886 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 177.483 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 147.820000 0.700000 148.200000 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.1284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.68 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 193.570000 200.100000 193.950000 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.9884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 191.130000 200.100000 191.510000 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 188.080000 200.100000 188.460000 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 185.030000 200.100000 185.410000 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 181.980000 200.100000 182.360000 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 179.540000 200.100000 179.920000 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 176.490000 200.100000 176.870000 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 173.440000 200.100000 173.820000 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 170.390000 200.100000 170.770000 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 167.340000 200.100000 167.720000 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 164.900000 200.100000 165.280000 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 161.850000 200.100000 162.230000 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 158.800000 200.100000 159.180000 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 155.750000 200.100000 156.130000 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.7824 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.168 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 153.310000 200.100000 153.690000 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.3684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.96 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 150.260000 200.100000 150.640000 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 147.210000 200.100000 147.590000 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 144.160000 200.100000 144.540000 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 141.110000 200.100000 141.490000 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 138.670000 200.100000 139.050000 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.4114 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.856 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 135.620000 200.100000 136.000000 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.7184 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.16 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 132.570000 200.100000 132.950000 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.2114 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.456 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 129.520000 200.100000 129.900000 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.9204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.904 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 126.470000 200.100000 126.850000 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.5214 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.776 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 124.030000 200.100000 124.410000 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.1324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.368 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 120.980000 200.100000 121.360000 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.648 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 117.930000 200.100000 118.310000 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.0624 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 114.880000 200.100000 115.260000 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.8884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.4 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 112.440000 200.100000 112.820000 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.5784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.08 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 109.390000 200.100000 109.770000 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.6144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.272 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 106.340000 200.100000 106.720000 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.5214 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.776 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 103.290000 200.100000 103.670000 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7103 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.3905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.3388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 140.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 57.7706 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 299.845 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 194.160000 0.000000 194.540000 0.700000 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.2798 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 96.173 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 33.2772 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 163.853 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 192.780000 0.000000 193.160000 0.700000 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.0422 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 89.985 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 26.995 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 133.435 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 191.400000 0.000000 191.780000 0.700000 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.2466 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 91.007 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 25.102 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 123.97 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 190.020000 0.000000 190.400000 0.700000 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.4062 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 91.805 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 27.8963 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 137.941 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 188.180000 0.000000 188.560000 0.700000 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.7115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.8888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 49.5801 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 257.434 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 186.800000 0.000000 187.180000 0.700000 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.9704 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 94.626 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 27.6702 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 135.52 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 185.420000 0.000000 185.800000 0.700000 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.2984 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 91.266 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 26.3634 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 130.277 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 183.580000 0.000000 183.960000 0.700000 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.3394 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 86.471 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 25.1444 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 123.486 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 182.200000 0.000000 182.580000 0.700000 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.6726 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 88.137 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 24.5024 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 120.972 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 180.820000 0.000000 181.200000 0.700000 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.1696 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 90.622 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 25.6054 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 126.487 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 179.440000 0.000000 179.820000 0.700000 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.4342 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 91.945 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 26.1182 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 129.051 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 177.600000 0.000000 177.980000 0.700000 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.0058 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 89.803 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 25.1246 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 124.083 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 176.220000 0.000000 176.600000 0.700000 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.5462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 92.505 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 25.4382 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 125.742 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 174.840000 0.000000 175.220000 0.700000 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.8322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 88.935 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 24.4766 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 120.934 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 173.000000 0.000000 173.380000 0.700000 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.7682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 83.615 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 25.3982 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 124.16 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 171.620000 0.000000 172.000000 0.700000 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.2918 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 86.233 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 24.8654 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 122.091 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 170.240000 0.000000 170.620000 0.700000 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.9652 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 89.6 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 24.6558 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 121.83 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 168.400000 0.000000 168.780000 0.700000 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8773 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.2255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.4788 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 163.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 60.8846 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 317.364 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 167.020000 0.000000 167.400000 0.700000 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.7098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.889 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3765 LAYER met2  ;
    ANTENNAMAXAREACAR 24.6455 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 114.047 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.46478 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 165.640000 0.000000 166.020000 0.700000 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.533 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.439 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 34.540000 199.560000 34.920000 200.260000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.249 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 32.700000 199.560000 33.080000 200.260000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.4542 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.045 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 31.320000 199.560000 31.700000 200.260000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.1252 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.4 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 29.940000 199.560000 30.320000 200.260000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.8874 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.329 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 28.560000 199.560000 28.940000 200.260000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.5186 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.367 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 27.180000 199.560000 27.560000 200.260000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.412 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 25.340000 199.560000 25.720000 200.260000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.0776 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.162 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 23.960000 199.560000 24.340000 200.260000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.0396 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.09 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 22.580000 199.560000 22.960000 200.260000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.8567 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.1225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.6148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.416 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 21.200000 199.560000 21.580000 200.260000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.009 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 19.360000 199.560000 19.740000 200.260000 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.757 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.559 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 17.980000 199.560000 18.360000 200.260000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.009 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 16.600000 199.560000 16.980000 200.260000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.7474 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.629 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 15.220000 199.560000 15.600000 200.260000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.411 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.947 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 13.840000 199.560000 14.220000 200.260000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.1726 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.755 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 12.460000 199.560000 12.840000 200.260000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6859 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.2685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.7468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.12 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 10.620000 199.560000 11.000000 200.260000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.233 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 9.240000 199.560000 9.620000 200.260000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.335 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.567 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 7.860000 199.560000 8.240000 200.260000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6304 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.034 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 6.480000 199.560000 6.860000 200.260000 ;
    END
  END FrameStrobe_O[0]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 198.900000 195.020000 200.100000 196.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 195.020000 1.200000 196.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.900000 2.850000 200.100000 4.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 1.200000 4.050000 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.070000 199.060000 197.270000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.070000 0.000000 197.270000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 199.060000 4.030000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 0.000000 4.030000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 200.100000 4.050000 ;
        RECT 0.000000 195.020000 200.100000 196.220000 ;
        RECT 2.830000 4.860000 4.030000 5.340000 ;
        RECT 2.830000 10.300000 4.030000 10.780000 ;
        RECT 7.060000 4.860000 8.260000 5.340000 ;
        RECT 7.060000 10.300000 8.260000 10.780000 ;
        RECT 2.830000 15.740000 4.030000 16.220000 ;
        RECT 7.060000 15.740000 8.260000 16.220000 ;
        RECT 2.830000 21.180000 4.030000 21.660000 ;
        RECT 7.060000 21.180000 8.260000 21.660000 ;
        RECT 2.830000 37.500000 4.030000 37.980000 ;
        RECT 7.060000 37.500000 8.260000 37.980000 ;
        RECT 2.830000 26.620000 4.030000 27.100000 ;
        RECT 7.060000 26.620000 8.260000 27.100000 ;
        RECT 2.830000 32.060000 4.030000 32.540000 ;
        RECT 7.060000 32.060000 8.260000 32.540000 ;
        RECT 2.830000 42.940000 4.030000 43.420000 ;
        RECT 7.060000 42.940000 8.260000 43.420000 ;
        RECT 2.830000 48.380000 4.030000 48.860000 ;
        RECT 7.060000 48.380000 8.260000 48.860000 ;
        RECT 52.060000 21.180000 53.260000 21.660000 ;
        RECT 52.060000 15.740000 53.260000 16.220000 ;
        RECT 52.060000 10.300000 53.260000 10.780000 ;
        RECT 52.060000 4.860000 53.260000 5.340000 ;
        RECT 97.060000 21.180000 98.260000 21.660000 ;
        RECT 97.060000 15.740000 98.260000 16.220000 ;
        RECT 97.060000 10.300000 98.260000 10.780000 ;
        RECT 97.060000 4.860000 98.260000 5.340000 ;
        RECT 52.060000 26.620000 53.260000 27.100000 ;
        RECT 52.060000 32.060000 53.260000 32.540000 ;
        RECT 52.060000 37.500000 53.260000 37.980000 ;
        RECT 52.060000 42.940000 53.260000 43.420000 ;
        RECT 52.060000 48.380000 53.260000 48.860000 ;
        RECT 97.060000 26.620000 98.260000 27.100000 ;
        RECT 97.060000 32.060000 98.260000 32.540000 ;
        RECT 97.060000 37.500000 98.260000 37.980000 ;
        RECT 97.060000 42.940000 98.260000 43.420000 ;
        RECT 97.060000 48.380000 98.260000 48.860000 ;
        RECT 2.830000 53.820000 4.030000 54.300000 ;
        RECT 7.060000 53.820000 8.260000 54.300000 ;
        RECT 2.830000 59.260000 4.030000 59.740000 ;
        RECT 7.060000 59.260000 8.260000 59.740000 ;
        RECT 2.830000 64.700000 4.030000 65.180000 ;
        RECT 7.060000 64.700000 8.260000 65.180000 ;
        RECT 2.830000 70.140000 4.030000 70.620000 ;
        RECT 7.060000 70.140000 8.260000 70.620000 ;
        RECT 7.060000 81.020000 8.260000 81.500000 ;
        RECT 2.830000 81.020000 4.030000 81.500000 ;
        RECT 2.830000 75.580000 4.030000 76.060000 ;
        RECT 7.060000 75.580000 8.260000 76.060000 ;
        RECT 2.830000 86.460000 4.030000 86.940000 ;
        RECT 7.060000 86.460000 8.260000 86.940000 ;
        RECT 2.830000 91.900000 4.030000 92.380000 ;
        RECT 7.060000 91.900000 8.260000 92.380000 ;
        RECT 2.830000 97.340000 4.030000 97.820000 ;
        RECT 7.060000 97.340000 8.260000 97.820000 ;
        RECT 52.060000 70.140000 53.260000 70.620000 ;
        RECT 52.060000 53.820000 53.260000 54.300000 ;
        RECT 52.060000 59.260000 53.260000 59.740000 ;
        RECT 52.060000 64.700000 53.260000 65.180000 ;
        RECT 97.060000 53.820000 98.260000 54.300000 ;
        RECT 97.060000 59.260000 98.260000 59.740000 ;
        RECT 97.060000 64.700000 98.260000 65.180000 ;
        RECT 97.060000 70.140000 98.260000 70.620000 ;
        RECT 52.060000 75.580000 53.260000 76.060000 ;
        RECT 52.060000 81.020000 53.260000 81.500000 ;
        RECT 52.060000 86.460000 53.260000 86.940000 ;
        RECT 52.060000 91.900000 53.260000 92.380000 ;
        RECT 52.060000 97.340000 53.260000 97.820000 ;
        RECT 97.060000 75.580000 98.260000 76.060000 ;
        RECT 97.060000 81.020000 98.260000 81.500000 ;
        RECT 97.060000 86.460000 98.260000 86.940000 ;
        RECT 97.060000 91.900000 98.260000 92.380000 ;
        RECT 97.060000 97.340000 98.260000 97.820000 ;
        RECT 142.060000 4.860000 143.260000 5.340000 ;
        RECT 142.060000 10.300000 143.260000 10.780000 ;
        RECT 142.060000 15.740000 143.260000 16.220000 ;
        RECT 142.060000 21.180000 143.260000 21.660000 ;
        RECT 142.060000 26.620000 143.260000 27.100000 ;
        RECT 142.060000 32.060000 143.260000 32.540000 ;
        RECT 142.060000 37.500000 143.260000 37.980000 ;
        RECT 142.060000 42.940000 143.260000 43.420000 ;
        RECT 142.060000 48.380000 143.260000 48.860000 ;
        RECT 196.070000 4.860000 197.270000 5.340000 ;
        RECT 196.070000 10.300000 197.270000 10.780000 ;
        RECT 187.060000 4.860000 188.260000 5.340000 ;
        RECT 187.060000 10.300000 188.260000 10.780000 ;
        RECT 187.060000 15.740000 188.260000 16.220000 ;
        RECT 187.060000 21.180000 188.260000 21.660000 ;
        RECT 196.070000 21.180000 197.270000 21.660000 ;
        RECT 196.070000 15.740000 197.270000 16.220000 ;
        RECT 196.070000 37.500000 197.270000 37.980000 ;
        RECT 187.060000 37.500000 188.260000 37.980000 ;
        RECT 196.070000 26.620000 197.270000 27.100000 ;
        RECT 196.070000 32.060000 197.270000 32.540000 ;
        RECT 187.060000 26.620000 188.260000 27.100000 ;
        RECT 187.060000 32.060000 188.260000 32.540000 ;
        RECT 196.070000 42.940000 197.270000 43.420000 ;
        RECT 196.070000 48.380000 197.270000 48.860000 ;
        RECT 187.060000 42.940000 188.260000 43.420000 ;
        RECT 187.060000 48.380000 188.260000 48.860000 ;
        RECT 142.060000 70.140000 143.260000 70.620000 ;
        RECT 142.060000 64.700000 143.260000 65.180000 ;
        RECT 142.060000 59.260000 143.260000 59.740000 ;
        RECT 142.060000 53.820000 143.260000 54.300000 ;
        RECT 142.060000 75.580000 143.260000 76.060000 ;
        RECT 142.060000 81.020000 143.260000 81.500000 ;
        RECT 142.060000 86.460000 143.260000 86.940000 ;
        RECT 142.060000 91.900000 143.260000 92.380000 ;
        RECT 142.060000 97.340000 143.260000 97.820000 ;
        RECT 187.060000 59.260000 188.260000 59.740000 ;
        RECT 187.060000 53.820000 188.260000 54.300000 ;
        RECT 196.070000 59.260000 197.270000 59.740000 ;
        RECT 196.070000 53.820000 197.270000 54.300000 ;
        RECT 196.070000 64.700000 197.270000 65.180000 ;
        RECT 196.070000 70.140000 197.270000 70.620000 ;
        RECT 187.060000 70.140000 188.260000 70.620000 ;
        RECT 187.060000 64.700000 188.260000 65.180000 ;
        RECT 187.060000 75.580000 188.260000 76.060000 ;
        RECT 187.060000 81.020000 188.260000 81.500000 ;
        RECT 187.060000 86.460000 188.260000 86.940000 ;
        RECT 196.070000 86.460000 197.270000 86.940000 ;
        RECT 196.070000 81.020000 197.270000 81.500000 ;
        RECT 196.070000 75.580000 197.270000 76.060000 ;
        RECT 196.070000 91.900000 197.270000 92.380000 ;
        RECT 196.070000 97.340000 197.270000 97.820000 ;
        RECT 187.060000 91.900000 188.260000 92.380000 ;
        RECT 187.060000 97.340000 188.260000 97.820000 ;
        RECT 2.830000 102.780000 4.030000 103.260000 ;
        RECT 7.060000 102.780000 8.260000 103.260000 ;
        RECT 2.830000 108.220000 4.030000 108.700000 ;
        RECT 7.060000 108.220000 8.260000 108.700000 ;
        RECT 2.830000 113.660000 4.030000 114.140000 ;
        RECT 7.060000 113.660000 8.260000 114.140000 ;
        RECT 2.830000 119.100000 4.030000 119.580000 ;
        RECT 2.830000 124.540000 4.030000 125.020000 ;
        RECT 7.060000 119.100000 8.260000 119.580000 ;
        RECT 7.060000 124.540000 8.260000 125.020000 ;
        RECT 2.830000 129.980000 4.030000 130.460000 ;
        RECT 7.060000 129.980000 8.260000 130.460000 ;
        RECT 2.830000 135.420000 4.030000 135.900000 ;
        RECT 7.060000 135.420000 8.260000 135.900000 ;
        RECT 2.830000 140.860000 4.030000 141.340000 ;
        RECT 7.060000 140.860000 8.260000 141.340000 ;
        RECT 2.830000 146.300000 4.030000 146.780000 ;
        RECT 7.060000 146.300000 8.260000 146.780000 ;
        RECT 52.060000 124.540000 53.260000 125.020000 ;
        RECT 52.060000 119.100000 53.260000 119.580000 ;
        RECT 52.060000 113.660000 53.260000 114.140000 ;
        RECT 52.060000 108.220000 53.260000 108.700000 ;
        RECT 52.060000 102.780000 53.260000 103.260000 ;
        RECT 97.060000 124.540000 98.260000 125.020000 ;
        RECT 97.060000 113.660000 98.260000 114.140000 ;
        RECT 97.060000 108.220000 98.260000 108.700000 ;
        RECT 97.060000 102.780000 98.260000 103.260000 ;
        RECT 97.060000 119.100000 98.260000 119.580000 ;
        RECT 52.060000 129.980000 53.260000 130.460000 ;
        RECT 52.060000 135.420000 53.260000 135.900000 ;
        RECT 52.060000 140.860000 53.260000 141.340000 ;
        RECT 52.060000 146.300000 53.260000 146.780000 ;
        RECT 97.060000 129.980000 98.260000 130.460000 ;
        RECT 97.060000 135.420000 98.260000 135.900000 ;
        RECT 97.060000 140.860000 98.260000 141.340000 ;
        RECT 97.060000 146.300000 98.260000 146.780000 ;
        RECT 2.830000 162.620000 4.030000 163.100000 ;
        RECT 7.060000 162.620000 8.260000 163.100000 ;
        RECT 2.830000 151.740000 4.030000 152.220000 ;
        RECT 7.060000 151.740000 8.260000 152.220000 ;
        RECT 2.830000 157.180000 4.030000 157.660000 ;
        RECT 7.060000 157.180000 8.260000 157.660000 ;
        RECT 2.830000 168.060000 4.030000 168.540000 ;
        RECT 7.060000 168.060000 8.260000 168.540000 ;
        RECT 2.830000 173.500000 4.030000 173.980000 ;
        RECT 7.060000 173.500000 8.260000 173.980000 ;
        RECT 2.830000 178.940000 4.030000 179.420000 ;
        RECT 7.060000 178.940000 8.260000 179.420000 ;
        RECT 7.060000 184.380000 8.260000 184.860000 ;
        RECT 2.830000 184.380000 4.030000 184.860000 ;
        RECT 2.830000 189.820000 4.030000 190.300000 ;
        RECT 7.060000 189.820000 8.260000 190.300000 ;
        RECT 52.060000 168.060000 53.260000 168.540000 ;
        RECT 52.060000 151.740000 53.260000 152.220000 ;
        RECT 52.060000 157.180000 53.260000 157.660000 ;
        RECT 52.060000 162.620000 53.260000 163.100000 ;
        RECT 52.060000 173.500000 53.260000 173.980000 ;
        RECT 97.060000 173.500000 98.260000 173.980000 ;
        RECT 97.060000 168.060000 98.260000 168.540000 ;
        RECT 97.060000 151.740000 98.260000 152.220000 ;
        RECT 97.060000 157.180000 98.260000 157.660000 ;
        RECT 97.060000 162.620000 98.260000 163.100000 ;
        RECT 52.060000 178.940000 53.260000 179.420000 ;
        RECT 52.060000 184.380000 53.260000 184.860000 ;
        RECT 52.060000 189.820000 53.260000 190.300000 ;
        RECT 97.060000 178.940000 98.260000 179.420000 ;
        RECT 97.060000 184.380000 98.260000 184.860000 ;
        RECT 97.060000 189.820000 98.260000 190.300000 ;
        RECT 142.060000 124.540000 143.260000 125.020000 ;
        RECT 142.060000 102.780000 143.260000 103.260000 ;
        RECT 142.060000 108.220000 143.260000 108.700000 ;
        RECT 142.060000 113.660000 143.260000 114.140000 ;
        RECT 142.060000 119.100000 143.260000 119.580000 ;
        RECT 142.060000 129.980000 143.260000 130.460000 ;
        RECT 142.060000 135.420000 143.260000 135.900000 ;
        RECT 142.060000 140.860000 143.260000 141.340000 ;
        RECT 142.060000 146.300000 143.260000 146.780000 ;
        RECT 196.070000 102.780000 197.270000 103.260000 ;
        RECT 196.070000 108.220000 197.270000 108.700000 ;
        RECT 187.060000 102.780000 188.260000 103.260000 ;
        RECT 187.060000 108.220000 188.260000 108.700000 ;
        RECT 187.060000 124.540000 188.260000 125.020000 ;
        RECT 187.060000 113.660000 188.260000 114.140000 ;
        RECT 187.060000 119.100000 188.260000 119.580000 ;
        RECT 196.070000 124.540000 197.270000 125.020000 ;
        RECT 196.070000 119.100000 197.270000 119.580000 ;
        RECT 196.070000 113.660000 197.270000 114.140000 ;
        RECT 196.070000 129.980000 197.270000 130.460000 ;
        RECT 196.070000 135.420000 197.270000 135.900000 ;
        RECT 187.060000 129.980000 188.260000 130.460000 ;
        RECT 187.060000 135.420000 188.260000 135.900000 ;
        RECT 187.060000 140.860000 188.260000 141.340000 ;
        RECT 187.060000 146.300000 188.260000 146.780000 ;
        RECT 196.070000 146.300000 197.270000 146.780000 ;
        RECT 196.070000 140.860000 197.270000 141.340000 ;
        RECT 142.060000 168.060000 143.260000 168.540000 ;
        RECT 142.060000 162.620000 143.260000 163.100000 ;
        RECT 142.060000 157.180000 143.260000 157.660000 ;
        RECT 142.060000 151.740000 143.260000 152.220000 ;
        RECT 142.060000 173.500000 143.260000 173.980000 ;
        RECT 142.060000 178.940000 143.260000 179.420000 ;
        RECT 142.060000 184.380000 143.260000 184.860000 ;
        RECT 142.060000 189.820000 143.260000 190.300000 ;
        RECT 196.070000 162.620000 197.270000 163.100000 ;
        RECT 187.060000 162.620000 188.260000 163.100000 ;
        RECT 196.070000 151.740000 197.270000 152.220000 ;
        RECT 196.070000 157.180000 197.270000 157.660000 ;
        RECT 187.060000 157.180000 188.260000 157.660000 ;
        RECT 187.060000 151.740000 188.260000 152.220000 ;
        RECT 196.070000 168.060000 197.270000 168.540000 ;
        RECT 196.070000 173.500000 197.270000 173.980000 ;
        RECT 187.060000 168.060000 188.260000 168.540000 ;
        RECT 187.060000 173.500000 188.260000 173.980000 ;
        RECT 187.060000 178.940000 188.260000 179.420000 ;
        RECT 187.060000 184.380000 188.260000 184.860000 ;
        RECT 196.070000 184.380000 197.270000 184.860000 ;
        RECT 196.070000 178.940000 197.270000 179.420000 ;
        RECT 196.070000 189.820000 197.270000 190.300000 ;
        RECT 187.060000 189.820000 188.260000 190.300000 ;
      LAYER met4 ;
        RECT 2.830000 0.000000 4.030000 200.260000 ;
        RECT 7.060000 2.850000 8.260000 196.220000 ;
        RECT 52.060000 2.850000 53.260000 196.220000 ;
        RECT 97.060000 2.850000 98.260000 196.220000 ;
        RECT 196.070000 0.000000 197.270000 200.260000 ;
        RECT 142.060000 2.850000 143.260000 196.220000 ;
        RECT 187.060000 2.850000 188.260000 196.220000 ;
    END
# end of P/G power stripe data as pin

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 198.900000 196.820000 200.100000 198.020000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 196.820000 1.200000 198.020000 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.900000 1.050000 200.100000 2.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 1.200000 2.250000 ;
    END
    PORT
      LAYER met4 ;
        RECT 197.870000 199.060000 199.070000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 197.870000 0.000000 199.070000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 199.060000 2.230000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 0.000000 2.230000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 200.100000 2.250000 ;
        RECT 0.000000 196.820000 200.100000 198.020000 ;
        RECT 4.895000 100.060000 6.260000 100.540000 ;
        RECT 1.030000 100.060000 2.230000 100.540000 ;
        RECT 95.060000 100.060000 96.260000 100.540000 ;
        RECT 50.060000 100.060000 51.260000 100.540000 ;
        RECT 197.870000 100.060000 199.070000 100.540000 ;
        RECT 185.060000 100.060000 186.260000 100.540000 ;
        RECT 140.060000 100.060000 141.260000 100.540000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 1.030000 7.580000 2.230000 8.060000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 1.030000 18.460000 2.230000 18.940000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 1.030000 13.020000 2.230000 13.500000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
        RECT 1.030000 23.900000 2.230000 24.380000 ;
        RECT 4.895000 29.340000 6.260000 29.820000 ;
        RECT 1.030000 29.340000 2.230000 29.820000 ;
        RECT 4.895000 34.780000 6.260000 35.260000 ;
        RECT 1.030000 34.780000 2.230000 35.260000 ;
        RECT 4.895000 40.220000 6.260000 40.700000 ;
        RECT 1.030000 40.220000 2.230000 40.700000 ;
        RECT 4.895000 45.660000 6.260000 46.140000 ;
        RECT 1.030000 45.660000 2.230000 46.140000 ;
        RECT 50.060000 23.900000 51.260000 24.380000 ;
        RECT 50.060000 18.460000 51.260000 18.940000 ;
        RECT 50.060000 13.020000 51.260000 13.500000 ;
        RECT 50.060000 7.580000 51.260000 8.060000 ;
        RECT 95.060000 23.900000 96.260000 24.380000 ;
        RECT 95.060000 18.460000 96.260000 18.940000 ;
        RECT 95.060000 13.020000 96.260000 13.500000 ;
        RECT 95.060000 7.580000 96.260000 8.060000 ;
        RECT 50.060000 45.660000 51.260000 46.140000 ;
        RECT 50.060000 40.220000 51.260000 40.700000 ;
        RECT 50.060000 34.780000 51.260000 35.260000 ;
        RECT 50.060000 29.340000 51.260000 29.820000 ;
        RECT 95.060000 45.660000 96.260000 46.140000 ;
        RECT 95.060000 40.220000 96.260000 40.700000 ;
        RECT 95.060000 34.780000 96.260000 35.260000 ;
        RECT 95.060000 29.340000 96.260000 29.820000 ;
        RECT 4.895000 51.100000 6.260000 51.580000 ;
        RECT 1.030000 51.100000 2.230000 51.580000 ;
        RECT 4.895000 61.980000 6.260000 62.460000 ;
        RECT 1.030000 61.980000 2.230000 62.460000 ;
        RECT 4.895000 56.540000 6.260000 57.020000 ;
        RECT 1.030000 56.540000 2.230000 57.020000 ;
        RECT 4.895000 67.420000 6.260000 67.900000 ;
        RECT 1.030000 67.420000 2.230000 67.900000 ;
        RECT 4.895000 72.860000 6.260000 73.340000 ;
        RECT 1.030000 72.860000 2.230000 73.340000 ;
        RECT 4.895000 78.300000 6.260000 78.780000 ;
        RECT 1.030000 78.300000 2.230000 78.780000 ;
        RECT 4.895000 83.740000 6.260000 84.220000 ;
        RECT 1.030000 83.740000 2.230000 84.220000 ;
        RECT 4.895000 89.180000 6.260000 89.660000 ;
        RECT 1.030000 89.180000 2.230000 89.660000 ;
        RECT 4.895000 94.620000 6.260000 95.100000 ;
        RECT 1.030000 94.620000 2.230000 95.100000 ;
        RECT 50.060000 72.860000 51.260000 73.340000 ;
        RECT 50.060000 67.420000 51.260000 67.900000 ;
        RECT 50.060000 61.980000 51.260000 62.460000 ;
        RECT 50.060000 56.540000 51.260000 57.020000 ;
        RECT 50.060000 51.100000 51.260000 51.580000 ;
        RECT 95.060000 72.860000 96.260000 73.340000 ;
        RECT 95.060000 67.420000 96.260000 67.900000 ;
        RECT 95.060000 61.980000 96.260000 62.460000 ;
        RECT 95.060000 56.540000 96.260000 57.020000 ;
        RECT 95.060000 51.100000 96.260000 51.580000 ;
        RECT 50.060000 94.620000 51.260000 95.100000 ;
        RECT 50.060000 89.180000 51.260000 89.660000 ;
        RECT 50.060000 83.740000 51.260000 84.220000 ;
        RECT 50.060000 78.300000 51.260000 78.780000 ;
        RECT 95.060000 94.620000 96.260000 95.100000 ;
        RECT 95.060000 89.180000 96.260000 89.660000 ;
        RECT 95.060000 83.740000 96.260000 84.220000 ;
        RECT 95.060000 78.300000 96.260000 78.780000 ;
        RECT 140.060000 23.900000 141.260000 24.380000 ;
        RECT 140.060000 18.460000 141.260000 18.940000 ;
        RECT 140.060000 13.020000 141.260000 13.500000 ;
        RECT 140.060000 7.580000 141.260000 8.060000 ;
        RECT 140.060000 45.660000 141.260000 46.140000 ;
        RECT 140.060000 40.220000 141.260000 40.700000 ;
        RECT 140.060000 34.780000 141.260000 35.260000 ;
        RECT 140.060000 29.340000 141.260000 29.820000 ;
        RECT 197.870000 7.580000 199.070000 8.060000 ;
        RECT 185.060000 7.580000 186.260000 8.060000 ;
        RECT 185.060000 13.020000 186.260000 13.500000 ;
        RECT 185.060000 18.460000 186.260000 18.940000 ;
        RECT 185.060000 23.900000 186.260000 24.380000 ;
        RECT 197.870000 23.900000 199.070000 24.380000 ;
        RECT 197.870000 13.020000 199.070000 13.500000 ;
        RECT 197.870000 18.460000 199.070000 18.940000 ;
        RECT 197.870000 34.780000 199.070000 35.260000 ;
        RECT 197.870000 29.340000 199.070000 29.820000 ;
        RECT 185.060000 34.780000 186.260000 35.260000 ;
        RECT 185.060000 29.340000 186.260000 29.820000 ;
        RECT 197.870000 45.660000 199.070000 46.140000 ;
        RECT 197.870000 40.220000 199.070000 40.700000 ;
        RECT 185.060000 45.660000 186.260000 46.140000 ;
        RECT 185.060000 40.220000 186.260000 40.700000 ;
        RECT 140.060000 72.860000 141.260000 73.340000 ;
        RECT 140.060000 67.420000 141.260000 67.900000 ;
        RECT 140.060000 61.980000 141.260000 62.460000 ;
        RECT 140.060000 56.540000 141.260000 57.020000 ;
        RECT 140.060000 51.100000 141.260000 51.580000 ;
        RECT 140.060000 94.620000 141.260000 95.100000 ;
        RECT 140.060000 89.180000 141.260000 89.660000 ;
        RECT 140.060000 83.740000 141.260000 84.220000 ;
        RECT 140.060000 78.300000 141.260000 78.780000 ;
        RECT 185.060000 51.100000 186.260000 51.580000 ;
        RECT 185.060000 56.540000 186.260000 57.020000 ;
        RECT 185.060000 61.980000 186.260000 62.460000 ;
        RECT 197.870000 61.980000 199.070000 62.460000 ;
        RECT 197.870000 51.100000 199.070000 51.580000 ;
        RECT 197.870000 56.540000 199.070000 57.020000 ;
        RECT 197.870000 72.860000 199.070000 73.340000 ;
        RECT 197.870000 67.420000 199.070000 67.900000 ;
        RECT 185.060000 72.860000 186.260000 73.340000 ;
        RECT 185.060000 67.420000 186.260000 67.900000 ;
        RECT 185.060000 78.300000 186.260000 78.780000 ;
        RECT 185.060000 83.740000 186.260000 84.220000 ;
        RECT 197.870000 83.740000 199.070000 84.220000 ;
        RECT 197.870000 78.300000 199.070000 78.780000 ;
        RECT 197.870000 94.620000 199.070000 95.100000 ;
        RECT 197.870000 89.180000 199.070000 89.660000 ;
        RECT 185.060000 94.620000 186.260000 95.100000 ;
        RECT 185.060000 89.180000 186.260000 89.660000 ;
        RECT 4.895000 105.500000 6.260000 105.980000 ;
        RECT 1.030000 105.500000 2.230000 105.980000 ;
        RECT 4.895000 110.940000 6.260000 111.420000 ;
        RECT 1.030000 110.940000 2.230000 111.420000 ;
        RECT 4.895000 116.380000 6.260000 116.860000 ;
        RECT 1.030000 116.380000 2.230000 116.860000 ;
        RECT 4.895000 121.820000 6.260000 122.300000 ;
        RECT 1.030000 121.820000 2.230000 122.300000 ;
        RECT 4.895000 127.260000 6.260000 127.740000 ;
        RECT 1.030000 127.260000 2.230000 127.740000 ;
        RECT 4.895000 132.700000 6.260000 133.180000 ;
        RECT 1.030000 132.700000 2.230000 133.180000 ;
        RECT 4.895000 143.580000 6.260000 144.060000 ;
        RECT 1.030000 143.580000 2.230000 144.060000 ;
        RECT 4.895000 138.140000 6.260000 138.620000 ;
        RECT 1.030000 138.140000 2.230000 138.620000 ;
        RECT 4.895000 149.020000 6.260000 149.500000 ;
        RECT 1.030000 149.020000 2.230000 149.500000 ;
        RECT 50.060000 121.820000 51.260000 122.300000 ;
        RECT 50.060000 116.380000 51.260000 116.860000 ;
        RECT 50.060000 110.940000 51.260000 111.420000 ;
        RECT 50.060000 105.500000 51.260000 105.980000 ;
        RECT 95.060000 121.820000 96.260000 122.300000 ;
        RECT 95.060000 116.380000 96.260000 116.860000 ;
        RECT 95.060000 110.940000 96.260000 111.420000 ;
        RECT 95.060000 105.500000 96.260000 105.980000 ;
        RECT 50.060000 149.020000 51.260000 149.500000 ;
        RECT 50.060000 143.580000 51.260000 144.060000 ;
        RECT 50.060000 138.140000 51.260000 138.620000 ;
        RECT 50.060000 132.700000 51.260000 133.180000 ;
        RECT 50.060000 127.260000 51.260000 127.740000 ;
        RECT 95.060000 149.020000 96.260000 149.500000 ;
        RECT 95.060000 143.580000 96.260000 144.060000 ;
        RECT 95.060000 138.140000 96.260000 138.620000 ;
        RECT 95.060000 132.700000 96.260000 133.180000 ;
        RECT 95.060000 127.260000 96.260000 127.740000 ;
        RECT 4.895000 154.460000 6.260000 154.940000 ;
        RECT 1.030000 154.460000 2.230000 154.940000 ;
        RECT 4.895000 159.900000 6.260000 160.380000 ;
        RECT 1.030000 159.900000 2.230000 160.380000 ;
        RECT 4.895000 165.340000 6.260000 165.820000 ;
        RECT 1.030000 165.340000 2.230000 165.820000 ;
        RECT 4.895000 170.780000 6.260000 171.260000 ;
        RECT 1.030000 170.780000 2.230000 171.260000 ;
        RECT 4.895000 176.220000 6.260000 176.700000 ;
        RECT 1.030000 176.220000 2.230000 176.700000 ;
        RECT 4.895000 187.100000 6.260000 187.580000 ;
        RECT 1.030000 187.100000 2.230000 187.580000 ;
        RECT 4.895000 181.660000 6.260000 182.140000 ;
        RECT 1.030000 181.660000 2.230000 182.140000 ;
        RECT 4.895000 192.540000 6.260000 193.020000 ;
        RECT 1.030000 192.540000 2.230000 193.020000 ;
        RECT 50.060000 170.780000 51.260000 171.260000 ;
        RECT 50.060000 165.340000 51.260000 165.820000 ;
        RECT 50.060000 159.900000 51.260000 160.380000 ;
        RECT 50.060000 154.460000 51.260000 154.940000 ;
        RECT 95.060000 170.780000 96.260000 171.260000 ;
        RECT 95.060000 165.340000 96.260000 165.820000 ;
        RECT 95.060000 159.900000 96.260000 160.380000 ;
        RECT 95.060000 154.460000 96.260000 154.940000 ;
        RECT 50.060000 192.540000 51.260000 193.020000 ;
        RECT 50.060000 187.100000 51.260000 187.580000 ;
        RECT 50.060000 181.660000 51.260000 182.140000 ;
        RECT 50.060000 176.220000 51.260000 176.700000 ;
        RECT 95.060000 192.540000 96.260000 193.020000 ;
        RECT 95.060000 187.100000 96.260000 187.580000 ;
        RECT 95.060000 176.220000 96.260000 176.700000 ;
        RECT 95.060000 181.660000 96.260000 182.140000 ;
        RECT 140.060000 121.820000 141.260000 122.300000 ;
        RECT 140.060000 116.380000 141.260000 116.860000 ;
        RECT 140.060000 110.940000 141.260000 111.420000 ;
        RECT 140.060000 105.500000 141.260000 105.980000 ;
        RECT 140.060000 149.020000 141.260000 149.500000 ;
        RECT 140.060000 143.580000 141.260000 144.060000 ;
        RECT 140.060000 138.140000 141.260000 138.620000 ;
        RECT 140.060000 132.700000 141.260000 133.180000 ;
        RECT 140.060000 127.260000 141.260000 127.740000 ;
        RECT 197.870000 110.940000 199.070000 111.420000 ;
        RECT 197.870000 105.500000 199.070000 105.980000 ;
        RECT 185.060000 110.940000 186.260000 111.420000 ;
        RECT 185.060000 105.500000 186.260000 105.980000 ;
        RECT 185.060000 116.380000 186.260000 116.860000 ;
        RECT 185.060000 121.820000 186.260000 122.300000 ;
        RECT 197.870000 121.820000 199.070000 122.300000 ;
        RECT 197.870000 116.380000 199.070000 116.860000 ;
        RECT 197.870000 132.700000 199.070000 133.180000 ;
        RECT 197.870000 127.260000 199.070000 127.740000 ;
        RECT 185.060000 132.700000 186.260000 133.180000 ;
        RECT 185.060000 127.260000 186.260000 127.740000 ;
        RECT 185.060000 138.140000 186.260000 138.620000 ;
        RECT 185.060000 143.580000 186.260000 144.060000 ;
        RECT 185.060000 149.020000 186.260000 149.500000 ;
        RECT 197.870000 149.020000 199.070000 149.500000 ;
        RECT 197.870000 138.140000 199.070000 138.620000 ;
        RECT 197.870000 143.580000 199.070000 144.060000 ;
        RECT 140.060000 170.780000 141.260000 171.260000 ;
        RECT 140.060000 165.340000 141.260000 165.820000 ;
        RECT 140.060000 154.460000 141.260000 154.940000 ;
        RECT 140.060000 159.900000 141.260000 160.380000 ;
        RECT 140.060000 192.540000 141.260000 193.020000 ;
        RECT 140.060000 187.100000 141.260000 187.580000 ;
        RECT 140.060000 181.660000 141.260000 182.140000 ;
        RECT 140.060000 176.220000 141.260000 176.700000 ;
        RECT 197.870000 159.900000 199.070000 160.380000 ;
        RECT 197.870000 154.460000 199.070000 154.940000 ;
        RECT 185.060000 159.900000 186.260000 160.380000 ;
        RECT 185.060000 154.460000 186.260000 154.940000 ;
        RECT 197.870000 170.780000 199.070000 171.260000 ;
        RECT 197.870000 165.340000 199.070000 165.820000 ;
        RECT 185.060000 170.780000 186.260000 171.260000 ;
        RECT 185.060000 165.340000 186.260000 165.820000 ;
        RECT 185.060000 176.220000 186.260000 176.700000 ;
        RECT 185.060000 181.660000 186.260000 182.140000 ;
        RECT 185.060000 187.100000 186.260000 187.580000 ;
        RECT 197.870000 187.100000 199.070000 187.580000 ;
        RECT 197.870000 176.220000 199.070000 176.700000 ;
        RECT 197.870000 181.660000 199.070000 182.140000 ;
        RECT 197.870000 192.540000 199.070000 193.020000 ;
        RECT 185.060000 192.540000 186.260000 193.020000 ;
      LAYER met4 ;
        RECT 1.030000 0.000000 2.230000 200.260000 ;
        RECT 5.060000 1.050000 6.260000 198.020000 ;
        RECT 50.060000 1.050000 51.260000 198.020000 ;
        RECT 95.060000 1.050000 96.260000 198.020000 ;
        RECT 197.870000 0.000000 199.070000 200.260000 ;
        RECT 140.060000 1.050000 141.260000 198.020000 ;
        RECT 185.060000 1.050000 186.260000 198.020000 ;
        RECT 4.895000 100.060000 6.260000 100.540000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
        RECT 4.895000 29.340000 6.260000 29.820000 ;
        RECT 4.895000 34.780000 6.260000 35.260000 ;
        RECT 4.895000 40.220000 6.260000 40.700000 ;
        RECT 4.895000 45.660000 6.260000 46.140000 ;
        RECT 4.895000 51.100000 6.260000 51.580000 ;
        RECT 4.895000 61.980000 6.260000 62.460000 ;
        RECT 4.895000 56.540000 6.260000 57.020000 ;
        RECT 4.895000 67.420000 6.260000 67.900000 ;
        RECT 4.895000 72.860000 6.260000 73.340000 ;
        RECT 4.895000 78.300000 6.260000 78.780000 ;
        RECT 4.895000 83.740000 6.260000 84.220000 ;
        RECT 4.895000 89.180000 6.260000 89.660000 ;
        RECT 4.895000 94.620000 6.260000 95.100000 ;
        RECT 4.895000 105.500000 6.260000 105.980000 ;
        RECT 4.895000 110.940000 6.260000 111.420000 ;
        RECT 4.895000 116.380000 6.260000 116.860000 ;
        RECT 4.895000 121.820000 6.260000 122.300000 ;
        RECT 4.895000 127.260000 6.260000 127.740000 ;
        RECT 4.895000 132.700000 6.260000 133.180000 ;
        RECT 4.895000 143.580000 6.260000 144.060000 ;
        RECT 4.895000 138.140000 6.260000 138.620000 ;
        RECT 4.895000 149.020000 6.260000 149.500000 ;
        RECT 4.895000 154.460000 6.260000 154.940000 ;
        RECT 4.895000 159.900000 6.260000 160.380000 ;
        RECT 4.895000 165.340000 6.260000 165.820000 ;
        RECT 4.895000 170.780000 6.260000 171.260000 ;
        RECT 4.895000 176.220000 6.260000 176.700000 ;
        RECT 4.895000 187.100000 6.260000 187.580000 ;
        RECT 4.895000 181.660000 6.260000 182.140000 ;
        RECT 4.895000 192.540000 6.260000 193.020000 ;
    END
# end of P/G power stripe data as pin

  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 200.100000 200.260000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 200.100000 200.260000 ;
    LAYER met2 ;
      RECT 35.060000 199.420000 200.100000 200.260000 ;
      RECT 33.220000 199.420000 34.400000 200.260000 ;
      RECT 31.840000 199.420000 32.560000 200.260000 ;
      RECT 30.460000 199.420000 31.180000 200.260000 ;
      RECT 29.080000 199.420000 29.800000 200.260000 ;
      RECT 27.700000 199.420000 28.420000 200.260000 ;
      RECT 25.860000 199.420000 27.040000 200.260000 ;
      RECT 24.480000 199.420000 25.200000 200.260000 ;
      RECT 23.100000 199.420000 23.820000 200.260000 ;
      RECT 21.720000 199.420000 22.440000 200.260000 ;
      RECT 19.880000 199.420000 21.060000 200.260000 ;
      RECT 18.500000 199.420000 19.220000 200.260000 ;
      RECT 17.120000 199.420000 17.840000 200.260000 ;
      RECT 15.740000 199.420000 16.460000 200.260000 ;
      RECT 14.360000 199.420000 15.080000 200.260000 ;
      RECT 12.980000 199.420000 13.700000 200.260000 ;
      RECT 11.140000 199.420000 12.320000 200.260000 ;
      RECT 9.760000 199.420000 10.480000 200.260000 ;
      RECT 8.380000 199.420000 9.100000 200.260000 ;
      RECT 7.000000 199.420000 7.720000 200.260000 ;
      RECT 5.620000 199.420000 6.340000 200.260000 ;
      RECT 0.000000 199.420000 4.960000 200.260000 ;
      RECT 0.000000 0.840000 200.100000 199.420000 ;
      RECT 194.680000 0.000000 200.100000 0.840000 ;
      RECT 193.300000 0.000000 194.020000 0.840000 ;
      RECT 191.920000 0.000000 192.640000 0.840000 ;
      RECT 190.540000 0.000000 191.260000 0.840000 ;
      RECT 188.700000 0.000000 189.880000 0.840000 ;
      RECT 187.320000 0.000000 188.040000 0.840000 ;
      RECT 185.940000 0.000000 186.660000 0.840000 ;
      RECT 184.100000 0.000000 185.280000 0.840000 ;
      RECT 182.720000 0.000000 183.440000 0.840000 ;
      RECT 181.340000 0.000000 182.060000 0.840000 ;
      RECT 179.960000 0.000000 180.680000 0.840000 ;
      RECT 178.120000 0.000000 179.300000 0.840000 ;
      RECT 176.740000 0.000000 177.460000 0.840000 ;
      RECT 175.360000 0.000000 176.080000 0.840000 ;
      RECT 173.520000 0.000000 174.700000 0.840000 ;
      RECT 172.140000 0.000000 172.860000 0.840000 ;
      RECT 170.760000 0.000000 171.480000 0.840000 ;
      RECT 168.920000 0.000000 170.100000 0.840000 ;
      RECT 167.540000 0.000000 168.260000 0.840000 ;
      RECT 166.160000 0.000000 166.880000 0.840000 ;
      RECT 164.780000 0.000000 165.500000 0.840000 ;
      RECT 162.940000 0.000000 164.120000 0.840000 ;
      RECT 161.560000 0.000000 162.280000 0.840000 ;
      RECT 160.180000 0.000000 160.900000 0.840000 ;
      RECT 158.340000 0.000000 159.520000 0.840000 ;
      RECT 156.960000 0.000000 157.680000 0.840000 ;
      RECT 155.580000 0.000000 156.300000 0.840000 ;
      RECT 154.200000 0.000000 154.920000 0.840000 ;
      RECT 152.360000 0.000000 153.540000 0.840000 ;
      RECT 150.980000 0.000000 151.700000 0.840000 ;
      RECT 149.600000 0.000000 150.320000 0.840000 ;
      RECT 147.760000 0.000000 148.940000 0.840000 ;
      RECT 146.380000 0.000000 147.100000 0.840000 ;
      RECT 145.000000 0.000000 145.720000 0.840000 ;
      RECT 143.160000 0.000000 144.340000 0.840000 ;
      RECT 141.780000 0.000000 142.500000 0.840000 ;
      RECT 140.400000 0.000000 141.120000 0.840000 ;
      RECT 139.020000 0.000000 139.740000 0.840000 ;
      RECT 137.180000 0.000000 138.360000 0.840000 ;
      RECT 135.800000 0.000000 136.520000 0.840000 ;
      RECT 134.420000 0.000000 135.140000 0.840000 ;
      RECT 132.580000 0.000000 133.760000 0.840000 ;
      RECT 131.200000 0.000000 131.920000 0.840000 ;
      RECT 129.820000 0.000000 130.540000 0.840000 ;
      RECT 127.980000 0.000000 129.160000 0.840000 ;
      RECT 126.600000 0.000000 127.320000 0.840000 ;
      RECT 125.220000 0.000000 125.940000 0.840000 ;
      RECT 123.840000 0.000000 124.560000 0.840000 ;
      RECT 122.000000 0.000000 123.180000 0.840000 ;
      RECT 120.620000 0.000000 121.340000 0.840000 ;
      RECT 119.240000 0.000000 119.960000 0.840000 ;
      RECT 117.400000 0.000000 118.580000 0.840000 ;
      RECT 116.020000 0.000000 116.740000 0.840000 ;
      RECT 114.640000 0.000000 115.360000 0.840000 ;
      RECT 113.260000 0.000000 113.980000 0.840000 ;
      RECT 111.420000 0.000000 112.600000 0.840000 ;
      RECT 110.040000 0.000000 110.760000 0.840000 ;
      RECT 108.660000 0.000000 109.380000 0.840000 ;
      RECT 106.820000 0.000000 108.000000 0.840000 ;
      RECT 105.440000 0.000000 106.160000 0.840000 ;
      RECT 104.060000 0.000000 104.780000 0.840000 ;
      RECT 102.220000 0.000000 103.400000 0.840000 ;
      RECT 100.840000 0.000000 101.560000 0.840000 ;
      RECT 99.460000 0.000000 100.180000 0.840000 ;
      RECT 98.080000 0.000000 98.800000 0.840000 ;
      RECT 96.240000 0.000000 97.420000 0.840000 ;
      RECT 94.860000 0.000000 95.580000 0.840000 ;
      RECT 93.480000 0.000000 94.200000 0.840000 ;
      RECT 91.640000 0.000000 92.820000 0.840000 ;
      RECT 90.260000 0.000000 90.980000 0.840000 ;
      RECT 88.880000 0.000000 89.600000 0.840000 ;
      RECT 87.040000 0.000000 88.220000 0.840000 ;
      RECT 85.660000 0.000000 86.380000 0.840000 ;
      RECT 84.280000 0.000000 85.000000 0.840000 ;
      RECT 82.900000 0.000000 83.620000 0.840000 ;
      RECT 81.060000 0.000000 82.240000 0.840000 ;
      RECT 79.680000 0.000000 80.400000 0.840000 ;
      RECT 78.300000 0.000000 79.020000 0.840000 ;
      RECT 76.460000 0.000000 77.640000 0.840000 ;
      RECT 75.080000 0.000000 75.800000 0.840000 ;
      RECT 73.700000 0.000000 74.420000 0.840000 ;
      RECT 72.320000 0.000000 73.040000 0.840000 ;
      RECT 70.480000 0.000000 71.660000 0.840000 ;
      RECT 69.100000 0.000000 69.820000 0.840000 ;
      RECT 67.720000 0.000000 68.440000 0.840000 ;
      RECT 65.880000 0.000000 67.060000 0.840000 ;
      RECT 64.500000 0.000000 65.220000 0.840000 ;
      RECT 63.120000 0.000000 63.840000 0.840000 ;
      RECT 61.280000 0.000000 62.460000 0.840000 ;
      RECT 59.900000 0.000000 60.620000 0.840000 ;
      RECT 58.520000 0.000000 59.240000 0.840000 ;
      RECT 57.140000 0.000000 57.860000 0.840000 ;
      RECT 55.300000 0.000000 56.480000 0.840000 ;
      RECT 53.920000 0.000000 54.640000 0.840000 ;
      RECT 52.540000 0.000000 53.260000 0.840000 ;
      RECT 50.700000 0.000000 51.880000 0.840000 ;
      RECT 49.320000 0.000000 50.040000 0.840000 ;
      RECT 47.940000 0.000000 48.660000 0.840000 ;
      RECT 46.100000 0.000000 47.280000 0.840000 ;
      RECT 44.720000 0.000000 45.440000 0.840000 ;
      RECT 43.340000 0.000000 44.060000 0.840000 ;
      RECT 41.960000 0.000000 42.680000 0.840000 ;
      RECT 40.120000 0.000000 41.300000 0.840000 ;
      RECT 38.740000 0.000000 39.460000 0.840000 ;
      RECT 37.360000 0.000000 38.080000 0.840000 ;
      RECT 35.520000 0.000000 36.700000 0.840000 ;
      RECT 34.140000 0.000000 34.860000 0.840000 ;
      RECT 32.760000 0.000000 33.480000 0.840000 ;
      RECT 31.380000 0.000000 32.100000 0.840000 ;
      RECT 29.540000 0.000000 30.720000 0.840000 ;
      RECT 28.160000 0.000000 28.880000 0.840000 ;
      RECT 26.780000 0.000000 27.500000 0.840000 ;
      RECT 24.940000 0.000000 26.120000 0.840000 ;
      RECT 23.560000 0.000000 24.280000 0.840000 ;
      RECT 22.180000 0.000000 22.900000 0.840000 ;
      RECT 20.340000 0.000000 21.520000 0.840000 ;
      RECT 18.960000 0.000000 19.680000 0.840000 ;
      RECT 17.580000 0.000000 18.300000 0.840000 ;
      RECT 16.200000 0.000000 16.920000 0.840000 ;
      RECT 14.360000 0.000000 15.540000 0.840000 ;
      RECT 12.980000 0.000000 13.700000 0.840000 ;
      RECT 11.600000 0.000000 12.320000 0.840000 ;
      RECT 9.760000 0.000000 10.940000 0.840000 ;
      RECT 8.380000 0.000000 9.100000 0.840000 ;
      RECT 7.000000 0.000000 7.720000 0.840000 ;
      RECT 5.620000 0.000000 6.340000 0.840000 ;
      RECT 0.000000 0.000000 4.960000 0.840000 ;
    LAYER met3 ;
      RECT 0.000000 198.320000 200.100000 200.260000 ;
      RECT 1.000000 194.250000 200.100000 194.720000 ;
      RECT 1.000000 193.880000 199.100000 194.250000 ;
      RECT 0.000000 193.320000 199.100000 193.880000 ;
      RECT 0.000000 193.030000 0.730000 193.320000 ;
      RECT 199.370000 192.240000 200.100000 193.270000 ;
      RECT 186.560000 192.240000 197.570000 193.320000 ;
      RECT 141.560000 192.240000 184.760000 193.320000 ;
      RECT 96.560000 192.240000 139.760000 193.320000 ;
      RECT 51.560000 192.240000 94.760000 193.320000 ;
      RECT 6.560000 192.240000 49.760000 193.320000 ;
      RECT 2.530000 192.240000 4.595000 193.320000 ;
      RECT 1.000000 192.050000 200.100000 192.240000 ;
      RECT 0.000000 191.810000 200.100000 192.050000 ;
      RECT 1.000000 190.830000 199.100000 191.810000 ;
      RECT 0.000000 190.600000 200.100000 190.830000 ;
      RECT 0.000000 189.980000 2.530000 190.600000 ;
      RECT 197.570000 189.520000 200.100000 190.600000 ;
      RECT 188.560000 189.520000 195.770000 190.600000 ;
      RECT 143.560000 189.520000 186.760000 190.600000 ;
      RECT 98.560000 189.520000 141.760000 190.600000 ;
      RECT 53.560000 189.520000 96.760000 190.600000 ;
      RECT 8.560000 189.520000 51.760000 190.600000 ;
      RECT 4.330000 189.520000 6.760000 190.600000 ;
      RECT 1.000000 189.520000 2.530000 189.980000 ;
      RECT 1.000000 189.000000 200.100000 189.520000 ;
      RECT 0.000000 188.760000 200.100000 189.000000 ;
      RECT 1.000000 187.880000 199.100000 188.760000 ;
      RECT 0.000000 186.930000 0.730000 187.780000 ;
      RECT 199.370000 186.800000 200.100000 187.780000 ;
      RECT 186.560000 186.800000 197.570000 187.880000 ;
      RECT 141.560000 186.800000 184.760000 187.880000 ;
      RECT 96.560000 186.800000 139.760000 187.880000 ;
      RECT 51.560000 186.800000 94.760000 187.880000 ;
      RECT 6.560000 186.800000 49.760000 187.880000 ;
      RECT 2.530000 186.800000 4.595000 187.880000 ;
      RECT 1.000000 185.950000 200.100000 186.800000 ;
      RECT 0.000000 185.710000 200.100000 185.950000 ;
      RECT 1.000000 185.160000 199.100000 185.710000 ;
      RECT 197.570000 184.730000 199.100000 185.160000 ;
      RECT 1.000000 184.730000 2.530000 185.160000 ;
      RECT 197.570000 184.080000 200.100000 184.730000 ;
      RECT 188.560000 184.080000 195.770000 185.160000 ;
      RECT 143.560000 184.080000 186.760000 185.160000 ;
      RECT 98.560000 184.080000 141.760000 185.160000 ;
      RECT 53.560000 184.080000 96.760000 185.160000 ;
      RECT 8.560000 184.080000 51.760000 185.160000 ;
      RECT 4.330000 184.080000 6.760000 185.160000 ;
      RECT 0.000000 184.080000 2.530000 184.730000 ;
      RECT 0.000000 183.880000 200.100000 184.080000 ;
      RECT 1.000000 182.900000 200.100000 183.880000 ;
      RECT 0.000000 182.660000 200.100000 182.900000 ;
      RECT 1.000000 182.440000 199.100000 182.660000 ;
      RECT 0.000000 181.440000 0.730000 181.680000 ;
      RECT 199.370000 181.360000 200.100000 181.680000 ;
      RECT 186.560000 181.360000 197.570000 182.440000 ;
      RECT 141.560000 181.360000 184.760000 182.440000 ;
      RECT 96.560000 181.360000 139.760000 182.440000 ;
      RECT 51.560000 181.360000 94.760000 182.440000 ;
      RECT 6.560000 181.360000 49.760000 182.440000 ;
      RECT 2.530000 181.360000 4.595000 182.440000 ;
      RECT 1.000000 180.460000 200.100000 181.360000 ;
      RECT 0.000000 180.220000 200.100000 180.460000 ;
      RECT 0.000000 179.720000 199.100000 180.220000 ;
      RECT 0.000000 179.610000 2.530000 179.720000 ;
      RECT 197.570000 179.240000 199.100000 179.720000 ;
      RECT 197.570000 178.640000 200.100000 179.240000 ;
      RECT 188.560000 178.640000 195.770000 179.720000 ;
      RECT 143.560000 178.640000 186.760000 179.720000 ;
      RECT 98.560000 178.640000 141.760000 179.720000 ;
      RECT 53.560000 178.640000 96.760000 179.720000 ;
      RECT 8.560000 178.640000 51.760000 179.720000 ;
      RECT 4.330000 178.640000 6.760000 179.720000 ;
      RECT 1.000000 178.640000 2.530000 179.610000 ;
      RECT 1.000000 178.630000 200.100000 178.640000 ;
      RECT 0.000000 178.390000 200.100000 178.630000 ;
      RECT 1.000000 177.410000 200.100000 178.390000 ;
      RECT 0.000000 177.170000 200.100000 177.410000 ;
      RECT 0.000000 177.000000 199.100000 177.170000 ;
      RECT 0.000000 176.560000 0.730000 177.000000 ;
      RECT 199.370000 175.920000 200.100000 176.190000 ;
      RECT 186.560000 175.920000 197.570000 177.000000 ;
      RECT 141.560000 175.920000 184.760000 177.000000 ;
      RECT 96.560000 175.920000 139.760000 177.000000 ;
      RECT 51.560000 175.920000 94.760000 177.000000 ;
      RECT 6.560000 175.920000 49.760000 177.000000 ;
      RECT 2.530000 175.920000 4.595000 177.000000 ;
      RECT 1.000000 175.580000 200.100000 175.920000 ;
      RECT 0.000000 175.340000 200.100000 175.580000 ;
      RECT 1.000000 174.360000 200.100000 175.340000 ;
      RECT 0.000000 174.280000 200.100000 174.360000 ;
      RECT 197.570000 174.120000 200.100000 174.280000 ;
      RECT 0.000000 173.510000 2.530000 174.280000 ;
      RECT 197.570000 173.200000 199.100000 174.120000 ;
      RECT 188.560000 173.200000 195.770000 174.280000 ;
      RECT 143.560000 173.200000 186.760000 174.280000 ;
      RECT 98.560000 173.200000 141.760000 174.280000 ;
      RECT 53.560000 173.200000 96.760000 174.280000 ;
      RECT 8.560000 173.200000 51.760000 174.280000 ;
      RECT 4.330000 173.200000 6.760000 174.280000 ;
      RECT 1.000000 173.200000 2.530000 173.510000 ;
      RECT 1.000000 173.140000 199.100000 173.200000 ;
      RECT 1.000000 172.530000 200.100000 173.140000 ;
      RECT 0.000000 172.290000 200.100000 172.530000 ;
      RECT 1.000000 171.560000 200.100000 172.290000 ;
      RECT 199.370000 171.070000 200.100000 171.560000 ;
      RECT 186.560000 170.480000 197.570000 171.560000 ;
      RECT 141.560000 170.480000 184.760000 171.560000 ;
      RECT 96.560000 170.480000 139.760000 171.560000 ;
      RECT 51.560000 170.480000 94.760000 171.560000 ;
      RECT 6.560000 170.480000 49.760000 171.560000 ;
      RECT 2.530000 170.480000 4.595000 171.560000 ;
      RECT 0.000000 170.480000 0.730000 171.310000 ;
      RECT 0.000000 170.460000 199.100000 170.480000 ;
      RECT 1.000000 170.090000 199.100000 170.460000 ;
      RECT 1.000000 169.480000 200.100000 170.090000 ;
      RECT 0.000000 169.240000 200.100000 169.480000 ;
      RECT 1.000000 168.840000 200.100000 169.240000 ;
      RECT 1.000000 168.260000 2.530000 168.840000 ;
      RECT 197.570000 168.020000 200.100000 168.840000 ;
      RECT 0.000000 168.020000 2.530000 168.260000 ;
      RECT 197.570000 167.760000 199.100000 168.020000 ;
      RECT 188.560000 167.760000 195.770000 168.840000 ;
      RECT 143.560000 167.760000 186.760000 168.840000 ;
      RECT 98.560000 167.760000 141.760000 168.840000 ;
      RECT 53.560000 167.760000 96.760000 168.840000 ;
      RECT 8.560000 167.760000 51.760000 168.840000 ;
      RECT 4.330000 167.760000 6.760000 168.840000 ;
      RECT 1.000000 167.760000 2.530000 168.020000 ;
      RECT 1.000000 167.040000 199.100000 167.760000 ;
      RECT 0.000000 166.190000 200.100000 167.040000 ;
      RECT 1.000000 166.120000 200.100000 166.190000 ;
      RECT 199.370000 165.580000 200.100000 166.120000 ;
      RECT 186.560000 165.040000 197.570000 166.120000 ;
      RECT 141.560000 165.040000 184.760000 166.120000 ;
      RECT 96.560000 165.040000 139.760000 166.120000 ;
      RECT 51.560000 165.040000 94.760000 166.120000 ;
      RECT 6.560000 165.040000 49.760000 166.120000 ;
      RECT 2.530000 165.040000 4.595000 166.120000 ;
      RECT 0.000000 165.040000 0.730000 165.210000 ;
      RECT 0.000000 164.970000 199.100000 165.040000 ;
      RECT 1.000000 164.600000 199.100000 164.970000 ;
      RECT 1.000000 163.990000 200.100000 164.600000 ;
      RECT 0.000000 163.400000 200.100000 163.990000 ;
      RECT 0.000000 163.140000 2.530000 163.400000 ;
      RECT 197.570000 162.530000 200.100000 163.400000 ;
      RECT 197.570000 162.320000 199.100000 162.530000 ;
      RECT 188.560000 162.320000 195.770000 163.400000 ;
      RECT 143.560000 162.320000 186.760000 163.400000 ;
      RECT 98.560000 162.320000 141.760000 163.400000 ;
      RECT 53.560000 162.320000 96.760000 163.400000 ;
      RECT 8.560000 162.320000 51.760000 163.400000 ;
      RECT 4.330000 162.320000 6.760000 163.400000 ;
      RECT 1.000000 162.320000 2.530000 163.140000 ;
      RECT 1.000000 162.160000 199.100000 162.320000 ;
      RECT 0.000000 161.920000 199.100000 162.160000 ;
      RECT 1.000000 161.550000 199.100000 161.920000 ;
      RECT 1.000000 160.940000 200.100000 161.550000 ;
      RECT 0.000000 160.680000 200.100000 160.940000 ;
      RECT 0.000000 160.090000 0.730000 160.680000 ;
      RECT 199.370000 159.600000 200.100000 160.680000 ;
      RECT 186.560000 159.600000 197.570000 160.680000 ;
      RECT 141.560000 159.600000 184.760000 160.680000 ;
      RECT 96.560000 159.600000 139.760000 160.680000 ;
      RECT 51.560000 159.600000 94.760000 160.680000 ;
      RECT 6.560000 159.600000 49.760000 160.680000 ;
      RECT 2.530000 159.600000 4.595000 160.680000 ;
      RECT 1.000000 159.480000 200.100000 159.600000 ;
      RECT 1.000000 159.110000 199.100000 159.480000 ;
      RECT 0.000000 158.870000 199.100000 159.110000 ;
      RECT 1.000000 158.500000 199.100000 158.870000 ;
      RECT 1.000000 157.960000 200.100000 158.500000 ;
      RECT 1.000000 157.890000 2.530000 157.960000 ;
      RECT 0.000000 157.040000 2.530000 157.890000 ;
      RECT 197.570000 156.880000 200.100000 157.960000 ;
      RECT 188.560000 156.880000 195.770000 157.960000 ;
      RECT 143.560000 156.880000 186.760000 157.960000 ;
      RECT 98.560000 156.880000 141.760000 157.960000 ;
      RECT 53.560000 156.880000 96.760000 157.960000 ;
      RECT 8.560000 156.880000 51.760000 157.960000 ;
      RECT 4.330000 156.880000 6.760000 157.960000 ;
      RECT 1.000000 156.880000 2.530000 157.040000 ;
      RECT 1.000000 156.430000 200.100000 156.880000 ;
      RECT 1.000000 156.060000 199.100000 156.430000 ;
      RECT 0.000000 155.820000 199.100000 156.060000 ;
      RECT 1.000000 155.450000 199.100000 155.820000 ;
      RECT 1.000000 155.240000 200.100000 155.450000 ;
      RECT 0.000000 154.600000 0.730000 154.840000 ;
      RECT 199.370000 154.160000 200.100000 155.240000 ;
      RECT 186.560000 154.160000 197.570000 155.240000 ;
      RECT 141.560000 154.160000 184.760000 155.240000 ;
      RECT 96.560000 154.160000 139.760000 155.240000 ;
      RECT 51.560000 154.160000 94.760000 155.240000 ;
      RECT 6.560000 154.160000 49.760000 155.240000 ;
      RECT 2.530000 154.160000 4.595000 155.240000 ;
      RECT 1.000000 153.990000 200.100000 154.160000 ;
      RECT 1.000000 153.620000 199.100000 153.990000 ;
      RECT 0.000000 153.010000 199.100000 153.620000 ;
      RECT 0.000000 152.770000 200.100000 153.010000 ;
      RECT 1.000000 152.520000 200.100000 152.770000 ;
      RECT 1.000000 151.790000 2.530000 152.520000 ;
      RECT 0.000000 151.550000 2.530000 151.790000 ;
      RECT 197.570000 151.440000 200.100000 152.520000 ;
      RECT 188.560000 151.440000 195.770000 152.520000 ;
      RECT 143.560000 151.440000 186.760000 152.520000 ;
      RECT 98.560000 151.440000 141.760000 152.520000 ;
      RECT 53.560000 151.440000 96.760000 152.520000 ;
      RECT 8.560000 151.440000 51.760000 152.520000 ;
      RECT 4.330000 151.440000 6.760000 152.520000 ;
      RECT 1.000000 151.440000 2.530000 151.550000 ;
      RECT 1.000000 150.940000 200.100000 151.440000 ;
      RECT 1.000000 150.570000 199.100000 150.940000 ;
      RECT 0.000000 149.960000 199.100000 150.570000 ;
      RECT 0.000000 149.800000 200.100000 149.960000 ;
      RECT 0.000000 149.720000 0.730000 149.800000 ;
      RECT 199.370000 148.720000 200.100000 149.800000 ;
      RECT 186.560000 148.720000 197.570000 149.800000 ;
      RECT 141.560000 148.720000 184.760000 149.800000 ;
      RECT 96.560000 148.720000 139.760000 149.800000 ;
      RECT 51.560000 148.720000 94.760000 149.800000 ;
      RECT 6.560000 148.720000 49.760000 149.800000 ;
      RECT 2.530000 148.720000 4.595000 149.800000 ;
      RECT 0.000000 148.720000 0.730000 148.740000 ;
      RECT 0.000000 148.500000 200.100000 148.720000 ;
      RECT 1.000000 147.890000 200.100000 148.500000 ;
      RECT 1.000000 147.520000 199.100000 147.890000 ;
      RECT 0.000000 147.080000 199.100000 147.520000 ;
      RECT 197.570000 146.910000 199.100000 147.080000 ;
      RECT 0.000000 146.670000 2.530000 147.080000 ;
      RECT 197.570000 146.000000 200.100000 146.910000 ;
      RECT 188.560000 146.000000 195.770000 147.080000 ;
      RECT 143.560000 146.000000 186.760000 147.080000 ;
      RECT 98.560000 146.000000 141.760000 147.080000 ;
      RECT 53.560000 146.000000 96.760000 147.080000 ;
      RECT 8.560000 146.000000 51.760000 147.080000 ;
      RECT 4.330000 146.000000 6.760000 147.080000 ;
      RECT 1.000000 146.000000 2.530000 146.670000 ;
      RECT 1.000000 145.690000 200.100000 146.000000 ;
      RECT 0.000000 145.450000 200.100000 145.690000 ;
      RECT 1.000000 144.840000 200.100000 145.450000 ;
      RECT 1.000000 144.470000 199.100000 144.840000 ;
      RECT 0.000000 144.360000 199.100000 144.470000 ;
      RECT 0.000000 144.230000 0.730000 144.360000 ;
      RECT 199.370000 143.280000 200.100000 143.860000 ;
      RECT 186.560000 143.280000 197.570000 144.360000 ;
      RECT 141.560000 143.280000 184.760000 144.360000 ;
      RECT 96.560000 143.280000 139.760000 144.360000 ;
      RECT 51.560000 143.280000 94.760000 144.360000 ;
      RECT 6.560000 143.280000 49.760000 144.360000 ;
      RECT 2.530000 143.280000 4.595000 144.360000 ;
      RECT 1.000000 143.250000 200.100000 143.280000 ;
      RECT 0.000000 142.400000 200.100000 143.250000 ;
      RECT 1.000000 141.790000 200.100000 142.400000 ;
      RECT 1.000000 141.640000 199.100000 141.790000 ;
      RECT 1.000000 141.420000 2.530000 141.640000 ;
      RECT 0.000000 141.180000 2.530000 141.420000 ;
      RECT 197.570000 140.810000 199.100000 141.640000 ;
      RECT 197.570000 140.560000 200.100000 140.810000 ;
      RECT 188.560000 140.560000 195.770000 141.640000 ;
      RECT 143.560000 140.560000 186.760000 141.640000 ;
      RECT 98.560000 140.560000 141.760000 141.640000 ;
      RECT 53.560000 140.560000 96.760000 141.640000 ;
      RECT 8.560000 140.560000 51.760000 141.640000 ;
      RECT 4.330000 140.560000 6.760000 141.640000 ;
      RECT 1.000000 140.560000 2.530000 141.180000 ;
      RECT 1.000000 140.200000 200.100000 140.560000 ;
      RECT 0.000000 139.350000 200.100000 140.200000 ;
      RECT 1.000000 138.920000 199.100000 139.350000 ;
      RECT 0.000000 138.130000 0.730000 138.370000 ;
      RECT 199.370000 137.840000 200.100000 138.370000 ;
      RECT 186.560000 137.840000 197.570000 138.920000 ;
      RECT 141.560000 137.840000 184.760000 138.920000 ;
      RECT 96.560000 137.840000 139.760000 138.920000 ;
      RECT 51.560000 137.840000 94.760000 138.920000 ;
      RECT 6.560000 137.840000 49.760000 138.920000 ;
      RECT 2.530000 137.840000 4.595000 138.920000 ;
      RECT 1.000000 137.150000 200.100000 137.840000 ;
      RECT 0.000000 136.300000 200.100000 137.150000 ;
      RECT 1.000000 136.200000 199.100000 136.300000 ;
      RECT 197.570000 135.320000 199.100000 136.200000 ;
      RECT 1.000000 135.320000 2.530000 136.200000 ;
      RECT 197.570000 135.120000 200.100000 135.320000 ;
      RECT 188.560000 135.120000 195.770000 136.200000 ;
      RECT 143.560000 135.120000 186.760000 136.200000 ;
      RECT 98.560000 135.120000 141.760000 136.200000 ;
      RECT 53.560000 135.120000 96.760000 136.200000 ;
      RECT 8.560000 135.120000 51.760000 136.200000 ;
      RECT 4.330000 135.120000 6.760000 136.200000 ;
      RECT 0.000000 135.120000 2.530000 135.320000 ;
      RECT 0.000000 135.080000 200.100000 135.120000 ;
      RECT 1.000000 134.100000 200.100000 135.080000 ;
      RECT 0.000000 133.480000 200.100000 134.100000 ;
      RECT 199.370000 133.250000 200.100000 133.480000 ;
      RECT 0.000000 133.250000 0.730000 133.480000 ;
      RECT 186.560000 132.400000 197.570000 133.480000 ;
      RECT 141.560000 132.400000 184.760000 133.480000 ;
      RECT 96.560000 132.400000 139.760000 133.480000 ;
      RECT 51.560000 132.400000 94.760000 133.480000 ;
      RECT 6.560000 132.400000 49.760000 133.480000 ;
      RECT 2.530000 132.400000 4.595000 133.480000 ;
      RECT 1.000000 132.270000 199.100000 132.400000 ;
      RECT 0.000000 132.030000 200.100000 132.270000 ;
      RECT 1.000000 131.050000 200.100000 132.030000 ;
      RECT 0.000000 130.810000 200.100000 131.050000 ;
      RECT 1.000000 130.760000 200.100000 130.810000 ;
      RECT 197.570000 130.200000 200.100000 130.760000 ;
      RECT 1.000000 129.830000 2.530000 130.760000 ;
      RECT 197.570000 129.680000 199.100000 130.200000 ;
      RECT 188.560000 129.680000 195.770000 130.760000 ;
      RECT 143.560000 129.680000 186.760000 130.760000 ;
      RECT 98.560000 129.680000 141.760000 130.760000 ;
      RECT 53.560000 129.680000 96.760000 130.760000 ;
      RECT 8.560000 129.680000 51.760000 130.760000 ;
      RECT 4.330000 129.680000 6.760000 130.760000 ;
      RECT 0.000000 129.680000 2.530000 129.830000 ;
      RECT 0.000000 129.220000 199.100000 129.680000 ;
      RECT 0.000000 128.980000 200.100000 129.220000 ;
      RECT 1.000000 128.040000 200.100000 128.980000 ;
      RECT 0.000000 127.760000 0.730000 128.000000 ;
      RECT 199.370000 127.150000 200.100000 128.040000 ;
      RECT 186.560000 126.960000 197.570000 128.040000 ;
      RECT 141.560000 126.960000 184.760000 128.040000 ;
      RECT 96.560000 126.960000 139.760000 128.040000 ;
      RECT 51.560000 126.960000 94.760000 128.040000 ;
      RECT 6.560000 126.960000 49.760000 128.040000 ;
      RECT 2.530000 126.960000 4.595000 128.040000 ;
      RECT 1.000000 126.780000 199.100000 126.960000 ;
      RECT 0.000000 126.170000 199.100000 126.780000 ;
      RECT 0.000000 125.930000 200.100000 126.170000 ;
      RECT 1.000000 125.320000 200.100000 125.930000 ;
      RECT 1.000000 124.950000 2.530000 125.320000 ;
      RECT 197.570000 124.710000 200.100000 125.320000 ;
      RECT 0.000000 124.710000 2.530000 124.950000 ;
      RECT 197.570000 124.240000 199.100000 124.710000 ;
      RECT 188.560000 124.240000 195.770000 125.320000 ;
      RECT 143.560000 124.240000 186.760000 125.320000 ;
      RECT 98.560000 124.240000 141.760000 125.320000 ;
      RECT 53.560000 124.240000 96.760000 125.320000 ;
      RECT 8.560000 124.240000 51.760000 125.320000 ;
      RECT 4.330000 124.240000 6.760000 125.320000 ;
      RECT 1.000000 124.240000 2.530000 124.710000 ;
      RECT 1.000000 123.730000 199.100000 124.240000 ;
      RECT 0.000000 122.880000 200.100000 123.730000 ;
      RECT 1.000000 122.600000 200.100000 122.880000 ;
      RECT 199.370000 121.660000 200.100000 122.600000 ;
      RECT 0.000000 121.660000 0.730000 121.900000 ;
      RECT 186.560000 121.520000 197.570000 122.600000 ;
      RECT 141.560000 121.520000 184.760000 122.600000 ;
      RECT 96.560000 121.520000 139.760000 122.600000 ;
      RECT 51.560000 121.520000 94.760000 122.600000 ;
      RECT 6.560000 121.520000 49.760000 122.600000 ;
      RECT 2.530000 121.520000 4.595000 122.600000 ;
      RECT 1.000000 120.680000 199.100000 121.520000 ;
      RECT 0.000000 119.880000 200.100000 120.680000 ;
      RECT 0.000000 119.830000 2.530000 119.880000 ;
      RECT 1.000000 118.850000 2.530000 119.830000 ;
      RECT 197.570000 118.800000 200.100000 119.880000 ;
      RECT 188.560000 118.800000 195.770000 119.880000 ;
      RECT 143.560000 118.800000 186.760000 119.880000 ;
      RECT 98.560000 118.800000 141.760000 119.880000 ;
      RECT 53.560000 118.800000 96.760000 119.880000 ;
      RECT 8.560000 118.800000 51.760000 119.880000 ;
      RECT 4.330000 118.800000 6.760000 119.880000 ;
      RECT 0.000000 118.800000 2.530000 118.850000 ;
      RECT 0.000000 118.610000 200.100000 118.800000 ;
      RECT 1.000000 117.630000 199.100000 118.610000 ;
      RECT 0.000000 117.390000 200.100000 117.630000 ;
      RECT 1.000000 117.160000 200.100000 117.390000 ;
      RECT 199.370000 116.080000 200.100000 117.160000 ;
      RECT 186.560000 116.080000 197.570000 117.160000 ;
      RECT 141.560000 116.080000 184.760000 117.160000 ;
      RECT 96.560000 116.080000 139.760000 117.160000 ;
      RECT 51.560000 116.080000 94.760000 117.160000 ;
      RECT 6.560000 116.080000 49.760000 117.160000 ;
      RECT 2.530000 116.080000 4.595000 117.160000 ;
      RECT 0.000000 116.080000 0.730000 116.410000 ;
      RECT 0.000000 115.560000 200.100000 116.080000 ;
      RECT 1.000000 114.580000 199.100000 115.560000 ;
      RECT 0.000000 114.440000 200.100000 114.580000 ;
      RECT 0.000000 114.340000 2.530000 114.440000 ;
      RECT 197.570000 113.360000 200.100000 114.440000 ;
      RECT 188.560000 113.360000 195.770000 114.440000 ;
      RECT 143.560000 113.360000 186.760000 114.440000 ;
      RECT 98.560000 113.360000 141.760000 114.440000 ;
      RECT 53.560000 113.360000 96.760000 114.440000 ;
      RECT 8.560000 113.360000 51.760000 114.440000 ;
      RECT 4.330000 113.360000 6.760000 114.440000 ;
      RECT 1.000000 113.360000 2.530000 114.340000 ;
      RECT 0.000000 113.120000 200.100000 113.360000 ;
      RECT 0.000000 112.510000 199.100000 113.120000 ;
      RECT 1.000000 112.140000 199.100000 112.510000 ;
      RECT 1.000000 111.720000 200.100000 112.140000 ;
      RECT 0.000000 111.290000 0.730000 111.530000 ;
      RECT 199.370000 110.640000 200.100000 111.720000 ;
      RECT 186.560000 110.640000 197.570000 111.720000 ;
      RECT 141.560000 110.640000 184.760000 111.720000 ;
      RECT 96.560000 110.640000 139.760000 111.720000 ;
      RECT 51.560000 110.640000 94.760000 111.720000 ;
      RECT 6.560000 110.640000 49.760000 111.720000 ;
      RECT 2.530000 110.640000 4.595000 111.720000 ;
      RECT 1.000000 110.310000 200.100000 110.640000 ;
      RECT 0.000000 110.070000 200.100000 110.310000 ;
      RECT 0.000000 109.460000 199.100000 110.070000 ;
      RECT 1.000000 109.090000 199.100000 109.460000 ;
      RECT 1.000000 109.000000 200.100000 109.090000 ;
      RECT 1.000000 108.480000 2.530000 109.000000 ;
      RECT 0.000000 108.240000 2.530000 108.480000 ;
      RECT 197.570000 107.920000 200.100000 109.000000 ;
      RECT 188.560000 107.920000 195.770000 109.000000 ;
      RECT 143.560000 107.920000 186.760000 109.000000 ;
      RECT 98.560000 107.920000 141.760000 109.000000 ;
      RECT 53.560000 107.920000 96.760000 109.000000 ;
      RECT 8.560000 107.920000 51.760000 109.000000 ;
      RECT 4.330000 107.920000 6.760000 109.000000 ;
      RECT 1.000000 107.920000 2.530000 108.240000 ;
      RECT 1.000000 107.260000 200.100000 107.920000 ;
      RECT 0.000000 107.020000 200.100000 107.260000 ;
      RECT 0.000000 106.410000 199.100000 107.020000 ;
      RECT 1.000000 106.280000 199.100000 106.410000 ;
      RECT 199.370000 105.200000 200.100000 106.040000 ;
      RECT 186.560000 105.200000 197.570000 106.280000 ;
      RECT 141.560000 105.200000 184.760000 106.280000 ;
      RECT 96.560000 105.200000 139.760000 106.280000 ;
      RECT 51.560000 105.200000 94.760000 106.280000 ;
      RECT 6.560000 105.200000 49.760000 106.280000 ;
      RECT 2.530000 105.200000 4.595000 106.280000 ;
      RECT 0.000000 105.200000 0.730000 105.430000 ;
      RECT 0.000000 105.190000 200.100000 105.200000 ;
      RECT 1.000000 104.210000 200.100000 105.190000 ;
      RECT 0.000000 103.970000 200.100000 104.210000 ;
      RECT 1.000000 103.560000 199.100000 103.970000 ;
      RECT 197.570000 102.990000 199.100000 103.560000 ;
      RECT 1.000000 102.990000 2.530000 103.560000 ;
      RECT 197.570000 102.480000 200.100000 102.990000 ;
      RECT 188.560000 102.480000 195.770000 103.560000 ;
      RECT 143.560000 102.480000 186.760000 103.560000 ;
      RECT 98.560000 102.480000 141.760000 103.560000 ;
      RECT 53.560000 102.480000 96.760000 103.560000 ;
      RECT 8.560000 102.480000 51.760000 103.560000 ;
      RECT 4.330000 102.480000 6.760000 103.560000 ;
      RECT 0.000000 102.480000 2.530000 102.990000 ;
      RECT 0.000000 102.140000 200.100000 102.480000 ;
      RECT 1.000000 101.160000 200.100000 102.140000 ;
      RECT 0.000000 100.920000 200.100000 101.160000 ;
      RECT 1.000000 100.840000 199.100000 100.920000 ;
      RECT 199.370000 99.760000 200.100000 99.940000 ;
      RECT 186.560000 99.760000 197.570000 100.840000 ;
      RECT 141.560000 99.760000 184.760000 100.840000 ;
      RECT 96.560000 99.760000 139.760000 100.840000 ;
      RECT 51.560000 99.760000 94.760000 100.840000 ;
      RECT 6.560000 99.760000 49.760000 100.840000 ;
      RECT 2.530000 99.760000 4.595000 100.840000 ;
      RECT 0.000000 99.760000 0.730000 99.940000 ;
      RECT 0.000000 99.090000 200.100000 99.760000 ;
      RECT 1.000000 98.480000 200.100000 99.090000 ;
      RECT 1.000000 98.120000 199.100000 98.480000 ;
      RECT 1.000000 98.110000 2.530000 98.120000 ;
      RECT 0.000000 97.870000 2.530000 98.110000 ;
      RECT 197.570000 97.500000 199.100000 98.120000 ;
      RECT 197.570000 97.040000 200.100000 97.500000 ;
      RECT 188.560000 97.040000 195.770000 98.120000 ;
      RECT 143.560000 97.040000 186.760000 98.120000 ;
      RECT 98.560000 97.040000 141.760000 98.120000 ;
      RECT 53.560000 97.040000 96.760000 98.120000 ;
      RECT 8.560000 97.040000 51.760000 98.120000 ;
      RECT 4.330000 97.040000 6.760000 98.120000 ;
      RECT 1.000000 97.040000 2.530000 97.870000 ;
      RECT 1.000000 96.890000 200.100000 97.040000 ;
      RECT 0.000000 96.040000 200.100000 96.890000 ;
      RECT 1.000000 95.430000 200.100000 96.040000 ;
      RECT 1.000000 95.400000 199.100000 95.430000 ;
      RECT 0.000000 94.820000 0.730000 95.060000 ;
      RECT 199.370000 94.320000 200.100000 94.450000 ;
      RECT 186.560000 94.320000 197.570000 95.400000 ;
      RECT 141.560000 94.320000 184.760000 95.400000 ;
      RECT 96.560000 94.320000 139.760000 95.400000 ;
      RECT 51.560000 94.320000 94.760000 95.400000 ;
      RECT 6.560000 94.320000 49.760000 95.400000 ;
      RECT 2.530000 94.320000 4.595000 95.400000 ;
      RECT 1.000000 93.840000 200.100000 94.320000 ;
      RECT 0.000000 93.600000 200.100000 93.840000 ;
      RECT 1.000000 92.680000 200.100000 93.600000 ;
      RECT 1.000000 92.620000 2.530000 92.680000 ;
      RECT 197.570000 92.380000 200.100000 92.680000 ;
      RECT 0.000000 91.770000 2.530000 92.620000 ;
      RECT 197.570000 91.600000 199.100000 92.380000 ;
      RECT 188.560000 91.600000 195.770000 92.680000 ;
      RECT 143.560000 91.600000 186.760000 92.680000 ;
      RECT 98.560000 91.600000 141.760000 92.680000 ;
      RECT 53.560000 91.600000 96.760000 92.680000 ;
      RECT 8.560000 91.600000 51.760000 92.680000 ;
      RECT 4.330000 91.600000 6.760000 92.680000 ;
      RECT 1.000000 91.600000 2.530000 91.770000 ;
      RECT 1.000000 91.400000 199.100000 91.600000 ;
      RECT 1.000000 90.790000 200.100000 91.400000 ;
      RECT 0.000000 90.550000 200.100000 90.790000 ;
      RECT 1.000000 89.960000 200.100000 90.550000 ;
      RECT 199.370000 89.330000 200.100000 89.960000 ;
      RECT 186.560000 88.880000 197.570000 89.960000 ;
      RECT 141.560000 88.880000 184.760000 89.960000 ;
      RECT 96.560000 88.880000 139.760000 89.960000 ;
      RECT 51.560000 88.880000 94.760000 89.960000 ;
      RECT 6.560000 88.880000 49.760000 89.960000 ;
      RECT 2.530000 88.880000 4.595000 89.960000 ;
      RECT 0.000000 88.880000 0.730000 89.570000 ;
      RECT 0.000000 88.720000 199.100000 88.880000 ;
      RECT 1.000000 88.350000 199.100000 88.720000 ;
      RECT 1.000000 87.740000 200.100000 88.350000 ;
      RECT 0.000000 87.500000 200.100000 87.740000 ;
      RECT 1.000000 87.240000 200.100000 87.500000 ;
      RECT 1.000000 86.520000 2.530000 87.240000 ;
      RECT 197.570000 86.280000 200.100000 87.240000 ;
      RECT 197.570000 86.160000 199.100000 86.280000 ;
      RECT 188.560000 86.160000 195.770000 87.240000 ;
      RECT 143.560000 86.160000 186.760000 87.240000 ;
      RECT 98.560000 86.160000 141.760000 87.240000 ;
      RECT 53.560000 86.160000 96.760000 87.240000 ;
      RECT 8.560000 86.160000 51.760000 87.240000 ;
      RECT 4.330000 86.160000 6.760000 87.240000 ;
      RECT 0.000000 86.160000 2.530000 86.520000 ;
      RECT 0.000000 85.670000 199.100000 86.160000 ;
      RECT 1.000000 85.300000 199.100000 85.670000 ;
      RECT 1.000000 84.690000 200.100000 85.300000 ;
      RECT 0.000000 84.520000 200.100000 84.690000 ;
      RECT 0.000000 84.450000 0.730000 84.520000 ;
      RECT 199.370000 83.840000 200.100000 84.520000 ;
      RECT 186.560000 83.440000 197.570000 84.520000 ;
      RECT 141.560000 83.440000 184.760000 84.520000 ;
      RECT 96.560000 83.440000 139.760000 84.520000 ;
      RECT 51.560000 83.440000 94.760000 84.520000 ;
      RECT 6.560000 83.440000 49.760000 84.520000 ;
      RECT 2.530000 83.440000 4.595000 84.520000 ;
      RECT 0.000000 83.440000 0.730000 83.470000 ;
      RECT 0.000000 82.860000 199.100000 83.440000 ;
      RECT 0.000000 82.620000 200.100000 82.860000 ;
      RECT 1.000000 81.800000 200.100000 82.620000 ;
      RECT 1.000000 81.640000 2.530000 81.800000 ;
      RECT 0.000000 81.400000 2.530000 81.640000 ;
      RECT 197.570000 80.790000 200.100000 81.800000 ;
      RECT 197.570000 80.720000 199.100000 80.790000 ;
      RECT 188.560000 80.720000 195.770000 81.800000 ;
      RECT 143.560000 80.720000 186.760000 81.800000 ;
      RECT 98.560000 80.720000 141.760000 81.800000 ;
      RECT 53.560000 80.720000 96.760000 81.800000 ;
      RECT 8.560000 80.720000 51.760000 81.800000 ;
      RECT 4.330000 80.720000 6.760000 81.800000 ;
      RECT 1.000000 80.720000 2.530000 81.400000 ;
      RECT 1.000000 80.420000 199.100000 80.720000 ;
      RECT 0.000000 80.180000 199.100000 80.420000 ;
      RECT 1.000000 79.810000 199.100000 80.180000 ;
      RECT 1.000000 79.200000 200.100000 79.810000 ;
      RECT 0.000000 79.080000 200.100000 79.200000 ;
      RECT 0.000000 78.350000 0.730000 79.080000 ;
      RECT 199.370000 78.000000 200.100000 79.080000 ;
      RECT 186.560000 78.000000 197.570000 79.080000 ;
      RECT 141.560000 78.000000 184.760000 79.080000 ;
      RECT 96.560000 78.000000 139.760000 79.080000 ;
      RECT 51.560000 78.000000 94.760000 79.080000 ;
      RECT 6.560000 78.000000 49.760000 79.080000 ;
      RECT 2.530000 78.000000 4.595000 79.080000 ;
      RECT 1.000000 77.740000 200.100000 78.000000 ;
      RECT 1.000000 77.370000 199.100000 77.740000 ;
      RECT 0.000000 77.130000 199.100000 77.370000 ;
      RECT 1.000000 76.760000 199.100000 77.130000 ;
      RECT 1.000000 76.360000 200.100000 76.760000 ;
      RECT 1.000000 76.150000 2.530000 76.360000 ;
      RECT 0.000000 75.300000 2.530000 76.150000 ;
      RECT 197.570000 75.280000 200.100000 76.360000 ;
      RECT 188.560000 75.280000 195.770000 76.360000 ;
      RECT 143.560000 75.280000 186.760000 76.360000 ;
      RECT 98.560000 75.280000 141.760000 76.360000 ;
      RECT 53.560000 75.280000 96.760000 76.360000 ;
      RECT 8.560000 75.280000 51.760000 76.360000 ;
      RECT 4.330000 75.280000 6.760000 76.360000 ;
      RECT 1.000000 75.280000 2.530000 75.300000 ;
      RECT 1.000000 74.690000 200.100000 75.280000 ;
      RECT 1.000000 74.320000 199.100000 74.690000 ;
      RECT 0.000000 74.080000 199.100000 74.320000 ;
      RECT 1.000000 73.710000 199.100000 74.080000 ;
      RECT 1.000000 73.640000 200.100000 73.710000 ;
      RECT 199.370000 72.560000 200.100000 73.640000 ;
      RECT 186.560000 72.560000 197.570000 73.640000 ;
      RECT 141.560000 72.560000 184.760000 73.640000 ;
      RECT 96.560000 72.560000 139.760000 73.640000 ;
      RECT 51.560000 72.560000 94.760000 73.640000 ;
      RECT 6.560000 72.560000 49.760000 73.640000 ;
      RECT 2.530000 72.560000 4.595000 73.640000 ;
      RECT 0.000000 72.560000 0.730000 73.100000 ;
      RECT 0.000000 72.250000 200.100000 72.560000 ;
      RECT 1.000000 71.270000 199.100000 72.250000 ;
      RECT 0.000000 71.030000 200.100000 71.270000 ;
      RECT 1.000000 70.920000 200.100000 71.030000 ;
      RECT 1.000000 70.050000 2.530000 70.920000 ;
      RECT 197.570000 69.840000 200.100000 70.920000 ;
      RECT 188.560000 69.840000 195.770000 70.920000 ;
      RECT 143.560000 69.840000 186.760000 70.920000 ;
      RECT 98.560000 69.840000 141.760000 70.920000 ;
      RECT 53.560000 69.840000 96.760000 70.920000 ;
      RECT 8.560000 69.840000 51.760000 70.920000 ;
      RECT 4.330000 69.840000 6.760000 70.920000 ;
      RECT 0.000000 69.840000 2.530000 70.050000 ;
      RECT 0.000000 69.200000 200.100000 69.840000 ;
      RECT 1.000000 68.220000 199.100000 69.200000 ;
      RECT 0.000000 68.200000 200.100000 68.220000 ;
      RECT 0.000000 67.980000 0.730000 68.200000 ;
      RECT 199.370000 67.120000 200.100000 68.200000 ;
      RECT 186.560000 67.120000 197.570000 68.200000 ;
      RECT 141.560000 67.120000 184.760000 68.200000 ;
      RECT 96.560000 67.120000 139.760000 68.200000 ;
      RECT 51.560000 67.120000 94.760000 68.200000 ;
      RECT 6.560000 67.120000 49.760000 68.200000 ;
      RECT 2.530000 67.120000 4.595000 68.200000 ;
      RECT 1.000000 67.000000 200.100000 67.120000 ;
      RECT 0.000000 66.760000 200.100000 67.000000 ;
      RECT 1.000000 66.150000 200.100000 66.760000 ;
      RECT 1.000000 65.780000 199.100000 66.150000 ;
      RECT 0.000000 65.480000 199.100000 65.780000 ;
      RECT 197.570000 65.170000 199.100000 65.480000 ;
      RECT 0.000000 64.930000 2.530000 65.480000 ;
      RECT 197.570000 64.400000 200.100000 65.170000 ;
      RECT 188.560000 64.400000 195.770000 65.480000 ;
      RECT 143.560000 64.400000 186.760000 65.480000 ;
      RECT 98.560000 64.400000 141.760000 65.480000 ;
      RECT 53.560000 64.400000 96.760000 65.480000 ;
      RECT 8.560000 64.400000 51.760000 65.480000 ;
      RECT 4.330000 64.400000 6.760000 65.480000 ;
      RECT 1.000000 64.400000 2.530000 64.930000 ;
      RECT 1.000000 63.950000 200.100000 64.400000 ;
      RECT 0.000000 63.710000 200.100000 63.950000 ;
      RECT 1.000000 63.100000 200.100000 63.710000 ;
      RECT 1.000000 62.760000 199.100000 63.100000 ;
      RECT 0.000000 61.880000 0.730000 62.730000 ;
      RECT 199.370000 61.680000 200.100000 62.120000 ;
      RECT 186.560000 61.680000 197.570000 62.760000 ;
      RECT 141.560000 61.680000 184.760000 62.760000 ;
      RECT 96.560000 61.680000 139.760000 62.760000 ;
      RECT 51.560000 61.680000 94.760000 62.760000 ;
      RECT 6.560000 61.680000 49.760000 62.760000 ;
      RECT 2.530000 61.680000 4.595000 62.760000 ;
      RECT 1.000000 60.900000 200.100000 61.680000 ;
      RECT 0.000000 60.660000 200.100000 60.900000 ;
      RECT 1.000000 60.050000 200.100000 60.660000 ;
      RECT 1.000000 60.040000 199.100000 60.050000 ;
      RECT 1.000000 59.680000 2.530000 60.040000 ;
      RECT 197.570000 59.070000 199.100000 60.040000 ;
      RECT 197.570000 58.960000 200.100000 59.070000 ;
      RECT 188.560000 58.960000 195.770000 60.040000 ;
      RECT 143.560000 58.960000 186.760000 60.040000 ;
      RECT 98.560000 58.960000 141.760000 60.040000 ;
      RECT 53.560000 58.960000 96.760000 60.040000 ;
      RECT 8.560000 58.960000 51.760000 60.040000 ;
      RECT 4.330000 58.960000 6.760000 60.040000 ;
      RECT 0.000000 58.960000 2.530000 59.680000 ;
      RECT 0.000000 58.830000 200.100000 58.960000 ;
      RECT 1.000000 57.850000 200.100000 58.830000 ;
      RECT 0.000000 57.610000 200.100000 57.850000 ;
      RECT 1.000000 57.320000 199.100000 57.610000 ;
      RECT 199.370000 56.240000 200.100000 56.630000 ;
      RECT 186.560000 56.240000 197.570000 57.320000 ;
      RECT 141.560000 56.240000 184.760000 57.320000 ;
      RECT 96.560000 56.240000 139.760000 57.320000 ;
      RECT 51.560000 56.240000 94.760000 57.320000 ;
      RECT 6.560000 56.240000 49.760000 57.320000 ;
      RECT 2.530000 56.240000 4.595000 57.320000 ;
      RECT 0.000000 56.240000 0.730000 56.630000 ;
      RECT 0.000000 55.780000 200.100000 56.240000 ;
      RECT 1.000000 54.800000 200.100000 55.780000 ;
      RECT 0.000000 54.600000 200.100000 54.800000 ;
      RECT 197.570000 54.560000 200.100000 54.600000 ;
      RECT 0.000000 54.560000 2.530000 54.600000 ;
      RECT 197.570000 53.580000 199.100000 54.560000 ;
      RECT 1.000000 53.580000 2.530000 54.560000 ;
      RECT 197.570000 53.520000 200.100000 53.580000 ;
      RECT 188.560000 53.520000 195.770000 54.600000 ;
      RECT 143.560000 53.520000 186.760000 54.600000 ;
      RECT 98.560000 53.520000 141.760000 54.600000 ;
      RECT 53.560000 53.520000 96.760000 54.600000 ;
      RECT 8.560000 53.520000 51.760000 54.600000 ;
      RECT 4.330000 53.520000 6.760000 54.600000 ;
      RECT 0.000000 53.520000 2.530000 53.580000 ;
      RECT 0.000000 53.340000 200.100000 53.520000 ;
      RECT 1.000000 52.360000 200.100000 53.340000 ;
      RECT 0.000000 51.880000 200.100000 52.360000 ;
      RECT 199.370000 51.510000 200.100000 51.880000 ;
      RECT 0.000000 51.510000 0.730000 51.880000 ;
      RECT 186.560000 50.800000 197.570000 51.880000 ;
      RECT 141.560000 50.800000 184.760000 51.880000 ;
      RECT 96.560000 50.800000 139.760000 51.880000 ;
      RECT 51.560000 50.800000 94.760000 51.880000 ;
      RECT 6.560000 50.800000 49.760000 51.880000 ;
      RECT 2.530000 50.800000 4.595000 51.880000 ;
      RECT 1.000000 50.530000 199.100000 50.800000 ;
      RECT 0.000000 50.290000 200.100000 50.530000 ;
      RECT 1.000000 49.310000 200.100000 50.290000 ;
      RECT 0.000000 49.160000 200.100000 49.310000 ;
      RECT 197.570000 48.460000 200.100000 49.160000 ;
      RECT 0.000000 48.460000 2.530000 49.160000 ;
      RECT 197.570000 48.080000 199.100000 48.460000 ;
      RECT 188.560000 48.080000 195.770000 49.160000 ;
      RECT 143.560000 48.080000 186.760000 49.160000 ;
      RECT 98.560000 48.080000 141.760000 49.160000 ;
      RECT 53.560000 48.080000 96.760000 49.160000 ;
      RECT 8.560000 48.080000 51.760000 49.160000 ;
      RECT 4.330000 48.080000 6.760000 49.160000 ;
      RECT 1.000000 48.080000 2.530000 48.460000 ;
      RECT 1.000000 47.480000 199.100000 48.080000 ;
      RECT 0.000000 47.240000 200.100000 47.480000 ;
      RECT 1.000000 46.440000 200.100000 47.240000 ;
      RECT 199.370000 46.020000 200.100000 46.440000 ;
      RECT 0.000000 45.410000 0.730000 46.260000 ;
      RECT 186.560000 45.360000 197.570000 46.440000 ;
      RECT 141.560000 45.360000 184.760000 46.440000 ;
      RECT 96.560000 45.360000 139.760000 46.440000 ;
      RECT 51.560000 45.360000 94.760000 46.440000 ;
      RECT 6.560000 45.360000 49.760000 46.440000 ;
      RECT 2.530000 45.360000 4.595000 46.440000 ;
      RECT 1.000000 45.040000 199.100000 45.360000 ;
      RECT 1.000000 44.430000 200.100000 45.040000 ;
      RECT 0.000000 44.190000 200.100000 44.430000 ;
      RECT 1.000000 43.720000 200.100000 44.190000 ;
      RECT 1.000000 43.210000 2.530000 43.720000 ;
      RECT 0.000000 42.970000 2.530000 43.210000 ;
      RECT 197.570000 42.640000 200.100000 43.720000 ;
      RECT 188.560000 42.640000 195.770000 43.720000 ;
      RECT 143.560000 42.640000 186.760000 43.720000 ;
      RECT 98.560000 42.640000 141.760000 43.720000 ;
      RECT 53.560000 42.640000 96.760000 43.720000 ;
      RECT 8.560000 42.640000 51.760000 43.720000 ;
      RECT 4.330000 42.640000 6.760000 43.720000 ;
      RECT 1.000000 42.640000 2.530000 42.970000 ;
      RECT 1.000000 41.990000 200.100000 42.640000 ;
      RECT 0.000000 41.140000 200.100000 41.990000 ;
      RECT 1.000000 41.000000 200.100000 41.140000 ;
      RECT 199.370000 39.920000 200.100000 41.000000 ;
      RECT 186.560000 39.920000 197.570000 41.000000 ;
      RECT 141.560000 39.920000 184.760000 41.000000 ;
      RECT 96.560000 39.920000 139.760000 41.000000 ;
      RECT 51.560000 39.920000 94.760000 41.000000 ;
      RECT 6.560000 39.920000 49.760000 41.000000 ;
      RECT 2.530000 39.920000 4.595000 41.000000 ;
      RECT 0.000000 39.920000 0.730000 40.160000 ;
      RECT 1.000000 38.940000 200.100000 39.920000 ;
      RECT 0.000000 38.280000 200.100000 38.940000 ;
      RECT 0.000000 38.090000 2.530000 38.280000 ;
      RECT 197.570000 37.200000 200.100000 38.280000 ;
      RECT 188.560000 37.200000 195.770000 38.280000 ;
      RECT 143.560000 37.200000 186.760000 38.280000 ;
      RECT 98.560000 37.200000 141.760000 38.280000 ;
      RECT 53.560000 37.200000 96.760000 38.280000 ;
      RECT 8.560000 37.200000 51.760000 38.280000 ;
      RECT 4.330000 37.200000 6.760000 38.280000 ;
      RECT 1.000000 37.200000 2.530000 38.090000 ;
      RECT 1.000000 37.110000 200.100000 37.200000 ;
      RECT 0.000000 36.870000 200.100000 37.110000 ;
      RECT 1.000000 35.890000 200.100000 36.870000 ;
      RECT 0.000000 35.560000 200.100000 35.890000 ;
      RECT 0.000000 35.040000 0.730000 35.560000 ;
      RECT 199.370000 34.480000 200.100000 35.560000 ;
      RECT 186.560000 34.480000 197.570000 35.560000 ;
      RECT 141.560000 34.480000 184.760000 35.560000 ;
      RECT 96.560000 34.480000 139.760000 35.560000 ;
      RECT 51.560000 34.480000 94.760000 35.560000 ;
      RECT 6.560000 34.480000 49.760000 35.560000 ;
      RECT 2.530000 34.480000 4.595000 35.560000 ;
      RECT 1.000000 34.060000 200.100000 34.480000 ;
      RECT 0.000000 33.820000 200.100000 34.060000 ;
      RECT 1.000000 32.840000 200.100000 33.820000 ;
      RECT 0.000000 31.990000 2.530000 32.840000 ;
      RECT 197.570000 31.760000 200.100000 32.840000 ;
      RECT 188.560000 31.760000 195.770000 32.840000 ;
      RECT 143.560000 31.760000 186.760000 32.840000 ;
      RECT 98.560000 31.760000 141.760000 32.840000 ;
      RECT 53.560000 31.760000 96.760000 32.840000 ;
      RECT 8.560000 31.760000 51.760000 32.840000 ;
      RECT 4.330000 31.760000 6.760000 32.840000 ;
      RECT 1.000000 31.760000 2.530000 31.990000 ;
      RECT 1.000000 31.010000 200.100000 31.760000 ;
      RECT 0.000000 30.770000 200.100000 31.010000 ;
      RECT 1.000000 30.120000 200.100000 30.770000 ;
      RECT 0.000000 29.550000 0.730000 29.790000 ;
      RECT 199.370000 29.040000 200.100000 30.120000 ;
      RECT 186.560000 29.040000 197.570000 30.120000 ;
      RECT 141.560000 29.040000 184.760000 30.120000 ;
      RECT 96.560000 29.040000 139.760000 30.120000 ;
      RECT 51.560000 29.040000 94.760000 30.120000 ;
      RECT 6.560000 29.040000 49.760000 30.120000 ;
      RECT 2.530000 29.040000 4.595000 30.120000 ;
      RECT 1.000000 28.570000 200.100000 29.040000 ;
      RECT 0.000000 27.720000 200.100000 28.570000 ;
      RECT 1.000000 27.400000 200.100000 27.720000 ;
      RECT 1.000000 26.740000 2.530000 27.400000 ;
      RECT 0.000000 26.500000 2.530000 26.740000 ;
      RECT 197.570000 26.320000 200.100000 27.400000 ;
      RECT 188.560000 26.320000 195.770000 27.400000 ;
      RECT 143.560000 26.320000 186.760000 27.400000 ;
      RECT 98.560000 26.320000 141.760000 27.400000 ;
      RECT 53.560000 26.320000 96.760000 27.400000 ;
      RECT 8.560000 26.320000 51.760000 27.400000 ;
      RECT 4.330000 26.320000 6.760000 27.400000 ;
      RECT 1.000000 26.320000 2.530000 26.500000 ;
      RECT 1.000000 25.520000 200.100000 26.320000 ;
      RECT 0.000000 24.680000 200.100000 25.520000 ;
      RECT 0.000000 24.670000 0.730000 24.680000 ;
      RECT 199.370000 23.600000 200.100000 24.680000 ;
      RECT 186.560000 23.600000 197.570000 24.680000 ;
      RECT 141.560000 23.600000 184.760000 24.680000 ;
      RECT 96.560000 23.600000 139.760000 24.680000 ;
      RECT 51.560000 23.600000 94.760000 24.680000 ;
      RECT 6.560000 23.600000 49.760000 24.680000 ;
      RECT 2.530000 23.600000 4.595000 24.680000 ;
      RECT 0.000000 23.600000 0.730000 23.690000 ;
      RECT 0.000000 23.450000 200.100000 23.600000 ;
      RECT 1.000000 22.470000 200.100000 23.450000 ;
      RECT 0.000000 21.960000 200.100000 22.470000 ;
      RECT 0.000000 21.620000 2.530000 21.960000 ;
      RECT 197.570000 20.880000 200.100000 21.960000 ;
      RECT 188.560000 20.880000 195.770000 21.960000 ;
      RECT 143.560000 20.880000 186.760000 21.960000 ;
      RECT 98.560000 20.880000 141.760000 21.960000 ;
      RECT 53.560000 20.880000 96.760000 21.960000 ;
      RECT 8.560000 20.880000 51.760000 21.960000 ;
      RECT 4.330000 20.880000 6.760000 21.960000 ;
      RECT 1.000000 20.880000 2.530000 21.620000 ;
      RECT 1.000000 20.640000 200.100000 20.880000 ;
      RECT 0.000000 20.400000 200.100000 20.640000 ;
      RECT 1.000000 19.420000 200.100000 20.400000 ;
      RECT 0.000000 19.240000 200.100000 19.420000 ;
      RECT 0.000000 18.570000 0.730000 19.240000 ;
      RECT 199.370000 18.160000 200.100000 19.240000 ;
      RECT 186.560000 18.160000 197.570000 19.240000 ;
      RECT 141.560000 18.160000 184.760000 19.240000 ;
      RECT 96.560000 18.160000 139.760000 19.240000 ;
      RECT 51.560000 18.160000 94.760000 19.240000 ;
      RECT 6.560000 18.160000 49.760000 19.240000 ;
      RECT 2.530000 18.160000 4.595000 19.240000 ;
      RECT 1.000000 17.590000 200.100000 18.160000 ;
      RECT 0.000000 17.350000 200.100000 17.590000 ;
      RECT 1.000000 16.520000 200.100000 17.350000 ;
      RECT 1.000000 16.370000 2.530000 16.520000 ;
      RECT 0.000000 16.130000 2.530000 16.370000 ;
      RECT 197.570000 15.440000 200.100000 16.520000 ;
      RECT 188.560000 15.440000 195.770000 16.520000 ;
      RECT 143.560000 15.440000 186.760000 16.520000 ;
      RECT 98.560000 15.440000 141.760000 16.520000 ;
      RECT 53.560000 15.440000 96.760000 16.520000 ;
      RECT 8.560000 15.440000 51.760000 16.520000 ;
      RECT 4.330000 15.440000 6.760000 16.520000 ;
      RECT 1.000000 15.440000 2.530000 16.130000 ;
      RECT 1.000000 15.150000 200.100000 15.440000 ;
      RECT 0.000000 14.300000 200.100000 15.150000 ;
      RECT 1.000000 13.800000 200.100000 14.300000 ;
      RECT 0.000000 13.080000 0.730000 13.320000 ;
      RECT 199.370000 12.720000 200.100000 13.800000 ;
      RECT 186.560000 12.720000 197.570000 13.800000 ;
      RECT 141.560000 12.720000 184.760000 13.800000 ;
      RECT 96.560000 12.720000 139.760000 13.800000 ;
      RECT 51.560000 12.720000 94.760000 13.800000 ;
      RECT 6.560000 12.720000 49.760000 13.800000 ;
      RECT 2.530000 12.720000 4.595000 13.800000 ;
      RECT 1.000000 12.100000 200.100000 12.720000 ;
      RECT 0.000000 11.250000 200.100000 12.100000 ;
      RECT 1.000000 11.080000 200.100000 11.250000 ;
      RECT 1.000000 10.270000 2.530000 11.080000 ;
      RECT 0.000000 10.030000 2.530000 10.270000 ;
      RECT 197.570000 10.000000 200.100000 11.080000 ;
      RECT 188.560000 10.000000 195.770000 11.080000 ;
      RECT 143.560000 10.000000 186.760000 11.080000 ;
      RECT 98.560000 10.000000 141.760000 11.080000 ;
      RECT 53.560000 10.000000 96.760000 11.080000 ;
      RECT 8.560000 10.000000 51.760000 11.080000 ;
      RECT 4.330000 10.000000 6.760000 11.080000 ;
      RECT 1.000000 10.000000 2.530000 10.030000 ;
      RECT 1.000000 9.050000 200.100000 10.000000 ;
      RECT 0.000000 8.360000 200.100000 9.050000 ;
      RECT 0.000000 8.200000 0.730000 8.360000 ;
      RECT 199.370000 7.280000 200.100000 8.360000 ;
      RECT 186.560000 7.280000 197.570000 8.360000 ;
      RECT 141.560000 7.280000 184.760000 8.360000 ;
      RECT 96.560000 7.280000 139.760000 8.360000 ;
      RECT 51.560000 7.280000 94.760000 8.360000 ;
      RECT 6.560000 7.280000 49.760000 8.360000 ;
      RECT 2.530000 7.280000 4.595000 8.360000 ;
      RECT 1.000000 7.220000 200.100000 7.280000 ;
      RECT 0.000000 6.980000 200.100000 7.220000 ;
      RECT 1.000000 6.000000 200.100000 6.980000 ;
      RECT 0.000000 5.760000 200.100000 6.000000 ;
      RECT 1.000000 5.640000 200.100000 5.760000 ;
      RECT 1.000000 4.780000 2.530000 5.640000 ;
      RECT 197.570000 4.560000 200.100000 5.640000 ;
      RECT 188.560000 4.560000 195.770000 5.640000 ;
      RECT 143.560000 4.560000 186.760000 5.640000 ;
      RECT 98.560000 4.560000 141.760000 5.640000 ;
      RECT 53.560000 4.560000 96.760000 5.640000 ;
      RECT 8.560000 4.560000 51.760000 5.640000 ;
      RECT 4.330000 4.560000 6.760000 5.640000 ;
      RECT 0.000000 4.560000 2.530000 4.780000 ;
      RECT 0.000000 4.350000 200.100000 4.560000 ;
      RECT 0.000000 0.000000 200.100000 0.750000 ;
    LAYER met4 ;
      RECT 4.330000 198.320000 195.770000 200.260000 ;
      RECT 186.560000 196.520000 195.770000 198.320000 ;
      RECT 141.560000 196.520000 184.760000 198.320000 ;
      RECT 96.560000 196.520000 139.760000 198.320000 ;
      RECT 51.560000 196.520000 94.760000 198.320000 ;
      RECT 6.560000 196.520000 49.760000 198.320000 ;
      RECT 4.330000 193.320000 4.760000 198.320000 ;
      RECT 4.330000 192.240000 4.595000 193.320000 ;
      RECT 4.330000 187.880000 4.760000 192.240000 ;
      RECT 4.330000 186.800000 4.595000 187.880000 ;
      RECT 4.330000 182.440000 4.760000 186.800000 ;
      RECT 4.330000 181.360000 4.595000 182.440000 ;
      RECT 4.330000 177.000000 4.760000 181.360000 ;
      RECT 4.330000 175.920000 4.595000 177.000000 ;
      RECT 4.330000 171.560000 4.760000 175.920000 ;
      RECT 4.330000 170.480000 4.595000 171.560000 ;
      RECT 4.330000 166.120000 4.760000 170.480000 ;
      RECT 4.330000 165.040000 4.595000 166.120000 ;
      RECT 4.330000 160.680000 4.760000 165.040000 ;
      RECT 4.330000 159.600000 4.595000 160.680000 ;
      RECT 4.330000 155.240000 4.760000 159.600000 ;
      RECT 4.330000 154.160000 4.595000 155.240000 ;
      RECT 4.330000 149.800000 4.760000 154.160000 ;
      RECT 4.330000 148.720000 4.595000 149.800000 ;
      RECT 4.330000 144.360000 4.760000 148.720000 ;
      RECT 4.330000 143.280000 4.595000 144.360000 ;
      RECT 4.330000 138.920000 4.760000 143.280000 ;
      RECT 4.330000 137.840000 4.595000 138.920000 ;
      RECT 4.330000 133.480000 4.760000 137.840000 ;
      RECT 4.330000 132.400000 4.595000 133.480000 ;
      RECT 4.330000 128.040000 4.760000 132.400000 ;
      RECT 4.330000 126.960000 4.595000 128.040000 ;
      RECT 4.330000 122.600000 4.760000 126.960000 ;
      RECT 4.330000 121.520000 4.595000 122.600000 ;
      RECT 4.330000 117.160000 4.760000 121.520000 ;
      RECT 4.330000 116.080000 4.595000 117.160000 ;
      RECT 4.330000 111.720000 4.760000 116.080000 ;
      RECT 4.330000 110.640000 4.595000 111.720000 ;
      RECT 4.330000 106.280000 4.760000 110.640000 ;
      RECT 4.330000 105.200000 4.595000 106.280000 ;
      RECT 4.330000 100.840000 4.760000 105.200000 ;
      RECT 4.330000 99.760000 4.595000 100.840000 ;
      RECT 4.330000 95.400000 4.760000 99.760000 ;
      RECT 4.330000 94.320000 4.595000 95.400000 ;
      RECT 4.330000 89.960000 4.760000 94.320000 ;
      RECT 4.330000 88.880000 4.595000 89.960000 ;
      RECT 4.330000 84.520000 4.760000 88.880000 ;
      RECT 4.330000 83.440000 4.595000 84.520000 ;
      RECT 4.330000 79.080000 4.760000 83.440000 ;
      RECT 4.330000 78.000000 4.595000 79.080000 ;
      RECT 4.330000 73.640000 4.760000 78.000000 ;
      RECT 4.330000 72.560000 4.595000 73.640000 ;
      RECT 4.330000 68.200000 4.760000 72.560000 ;
      RECT 4.330000 67.120000 4.595000 68.200000 ;
      RECT 4.330000 62.760000 4.760000 67.120000 ;
      RECT 4.330000 61.680000 4.595000 62.760000 ;
      RECT 4.330000 57.320000 4.760000 61.680000 ;
      RECT 4.330000 56.240000 4.595000 57.320000 ;
      RECT 4.330000 51.880000 4.760000 56.240000 ;
      RECT 4.330000 50.800000 4.595000 51.880000 ;
      RECT 4.330000 46.440000 4.760000 50.800000 ;
      RECT 4.330000 45.360000 4.595000 46.440000 ;
      RECT 4.330000 41.000000 4.760000 45.360000 ;
      RECT 4.330000 39.920000 4.595000 41.000000 ;
      RECT 4.330000 35.560000 4.760000 39.920000 ;
      RECT 4.330000 34.480000 4.595000 35.560000 ;
      RECT 4.330000 30.120000 4.760000 34.480000 ;
      RECT 4.330000 29.040000 4.595000 30.120000 ;
      RECT 4.330000 24.680000 4.760000 29.040000 ;
      RECT 4.330000 23.600000 4.595000 24.680000 ;
      RECT 4.330000 19.240000 4.760000 23.600000 ;
      RECT 4.330000 18.160000 4.595000 19.240000 ;
      RECT 4.330000 13.800000 4.760000 18.160000 ;
      RECT 4.330000 12.720000 4.595000 13.800000 ;
      RECT 4.330000 8.360000 4.760000 12.720000 ;
      RECT 4.330000 7.280000 4.595000 8.360000 ;
      RECT 188.560000 2.550000 195.770000 196.520000 ;
      RECT 186.560000 2.550000 186.760000 196.520000 ;
      RECT 143.560000 2.550000 184.760000 196.520000 ;
      RECT 141.560000 2.550000 141.760000 196.520000 ;
      RECT 98.560000 2.550000 139.760000 196.520000 ;
      RECT 96.560000 2.550000 96.760000 196.520000 ;
      RECT 53.560000 2.550000 94.760000 196.520000 ;
      RECT 51.560000 2.550000 51.760000 196.520000 ;
      RECT 8.560000 2.550000 49.760000 196.520000 ;
      RECT 6.560000 2.550000 6.760000 196.520000 ;
      RECT 186.560000 0.750000 195.770000 2.550000 ;
      RECT 141.560000 0.750000 184.760000 2.550000 ;
      RECT 96.560000 0.750000 139.760000 2.550000 ;
      RECT 51.560000 0.750000 94.760000 2.550000 ;
      RECT 6.560000 0.750000 49.760000 2.550000 ;
      RECT 4.330000 0.750000 4.760000 7.280000 ;
      RECT 199.370000 0.000000 200.100000 200.260000 ;
      RECT 4.330000 0.000000 195.770000 0.750000 ;
      RECT 0.000000 0.000000 0.730000 200.260000 ;
  END
END E_CPU_IO_bot

END LIBRARY
