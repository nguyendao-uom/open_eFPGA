##
## LEF for PtnCells ;
## created by Innovus v19.11-s128_1 on Thu Dec 23 11:01:41 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO flexbex_ibex_core
  CLASS BLOCK ;
  SIZE 550.160000 BY 549.780000 ;
  FOREIGN flexbex_ibex_core 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.2228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.992 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.608 LAYER met3  ;
    ANTENNAMAXAREACAR 1.52077 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 6.9847 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.0386502 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 10.160000 0.000000 10.540000 0.900000 ;
    END
  END clk_i
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5785 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4095 LAYER met2  ;
    ANTENNAMAXAREACAR 20.8916 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 98.763 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.354644 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4095 LAYER met3  ;
    ANTENNAMAXAREACAR 21.5143 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 103.178 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.452324 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 199.318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1066.77 LAYER met4  ;
    ANTENNAGATEAREA 3.087 LAYER met4  ;
    ANTENNAMAXAREACAR 135.617 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 721.122 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.804695 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 12.000000 0.000000 12.380000 0.900000 ;
    END
  END rst_ni
  PIN test_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.675 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.267 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 23.7444 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 109.679 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 14.300000 0.000000 14.680000 0.900000 ;
    END
  END test_en_i
  PIN core_id_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6121 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.2388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 135.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 63.8632 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 328.376 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 16.600000 0.000000 16.980000 0.900000 ;
    END
  END core_id_i[3]
  PIN core_id_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9927 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.5556 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 121.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.5588 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.784 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 34.5933 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 177.265 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 18.900000 0.000000 19.280000 0.900000 ;
    END
  END core_id_i[2]
  PIN core_id_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7093 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.1495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.5462 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 95.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.1838 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 54.784 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 50.0984 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 266.154 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 21.200000 0.000000 21.580000 0.900000 ;
    END
  END core_id_i[1]
  PIN core_id_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4413 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.4614 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 169.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.6698 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 41.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 40.2309 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 215.616 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 23.500000 0.000000 23.880000 0.900000 ;
    END
  END core_id_i[0]
  PIN cluster_id_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.1667 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 90.4365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.2628 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.872 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 54.744 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 288.012 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 25.800000 0.000000 26.180000 0.900000 ;
    END
  END cluster_id_i[5]
  PIN cluster_id_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0875 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.0405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.032 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 44.0838 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 224.764 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 28.100000 0.000000 28.480000 0.900000 ;
    END
  END cluster_id_i[4]
  PIN cluster_id_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2063 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.8605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.9968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 128.92 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.6504 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.88 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 22.1467 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 119.887 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 30.400000 0.000000 30.780000 0.900000 ;
    END
  END cluster_id_i[3]
  PIN cluster_id_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8613 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.8995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.1054 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.7666 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 63.696 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 62.6006 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 334.687 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 32.700000 0.000000 33.080000 0.900000 ;
    END
  END cluster_id_i[2]
  PIN cluster_id_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6963 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.9166 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.4336 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 21.1867 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 112.303 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 35.000000 0.000000 35.380000 0.900000 ;
    END
  END cluster_id_i[1]
  PIN cluster_id_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8683 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.6206 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 145.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 21.9016 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 117.701 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 37.300000 0.000000 37.680000 0.900000 ;
    END
  END cluster_id_i[0]
  PIN boot_addr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9327 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 28.3086 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 151.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 62.1553 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 325.181 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.423165 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 39.600000 0.000000 39.980000 0.900000 ;
    END
  END boot_addr_i[31]
  PIN boot_addr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1545 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.6115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 25.8348 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 138.256 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 54.205 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 280.343 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.423165 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 41.900000 0.000000 42.280000 0.900000 ;
    END
  END boot_addr_i[30]
  PIN boot_addr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2323 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.3855 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 242.992 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 84.923 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 445.196 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 44.200000 0.000000 44.580000 0.900000 ;
    END
  END boot_addr_i[29]
  PIN boot_addr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.2063 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.6345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.7174 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.904 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met3  ;
    ANTENNAMAXAREACAR 133.267 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 660.588 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 46.500000 0.000000 46.880000 0.900000 ;
    END
  END boot_addr_i[28]
  PIN boot_addr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.8853 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.2655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.8988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.1205 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 102.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 49.6966 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 255.696 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 48.800000 0.000000 49.180000 0.900000 ;
    END
  END boot_addr_i[27]
  PIN boot_addr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.4055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.2647 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 220.544 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 88.7349 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 462.746 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 51.100000 0.000000 51.480000 0.900000 ;
    END
  END boot_addr_i[26]
  PIN boot_addr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3821 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 44.1447 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 235.904 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 81.3654 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 426.703 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 53.400000 0.000000 53.780000 0.900000 ;
    END
  END boot_addr_i[25]
  PIN boot_addr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1401 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.125 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 40.5327 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 216.64 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 75.3498 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 393.785 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 55.700000 0.000000 56.080000 0.900000 ;
    END
  END boot_addr_i[24]
  PIN boot_addr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4305 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.791 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.5917 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 222.288 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 87.921 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 460.666 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 58.000000 0.000000 58.380000 0.900000 ;
    END
  END boot_addr_i[23]
  PIN boot_addr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.885 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 37.8267 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 202.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 67.9423 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 355.117 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 60.300000 0.000000 60.680000 0.900000 ;
    END
  END boot_addr_i[22]
  PIN boot_addr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4489 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.0835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.8565 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 181.504 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 65.4832 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 341.61 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 62.600000 0.000000 62.980000 0.900000 ;
    END
  END boot_addr_i[21]
  PIN boot_addr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7089 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.3835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.645 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.0297 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 176.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 61.3685 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 320.204 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 64.900000 0.000000 65.280000 0.900000 ;
    END
  END boot_addr_i[20]
  PIN boot_addr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7103 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.3905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.713 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.4087 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 157.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 65.5137 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 339.535 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 67.200000 0.000000 67.580000 0.900000 ;
    END
  END boot_addr_i[19]
  PIN boot_addr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.689 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 40.8747 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 218.464 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 76.537 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 400.088 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 69.500000 0.000000 69.880000 0.900000 ;
    END
  END boot_addr_i[18]
  PIN boot_addr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4183 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.9305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.896 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.8337 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 148.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 55.2712 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 287.111 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 71.800000 0.000000 72.180000 0.900000 ;
    END
  END boot_addr_i[17]
  PIN boot_addr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 40.1187 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 214.432 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 94.6347 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 495.817 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 74.100000 0.000000 74.480000 0.900000 ;
    END
  END boot_addr_i[16]
  PIN boot_addr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.5107 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 221.856 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 73.0112 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 386.006 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 76.400000 0.000000 76.780000 0.900000 ;
    END
  END boot_addr_i[15]
  PIN boot_addr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2533 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.1055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.492 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 39.3957 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 210.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 79.2864 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 415.766 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 78.700000 0.000000 79.080000 0.900000 ;
    END
  END boot_addr_i[14]
  PIN boot_addr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 37.3737 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 199.792 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 86.1787 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 447.147 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 81.000000 0.000000 81.380000 0.900000 ;
    END
  END boot_addr_i[13]
  PIN boot_addr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8683 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.6876 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 180.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 52.1101 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 275.166 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 83.300000 0.000000 83.680000 0.900000 ;
    END
  END boot_addr_i[12]
  PIN boot_addr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.5928 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 147.632 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 46.9526 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 244.925 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.315421 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 85.600000 0.000000 85.980000 0.900000 ;
    END
  END boot_addr_i[11]
  PIN boot_addr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 40.5327 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 216.64 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 61.0485 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 322.781 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 87.900000 0.000000 88.280000 0.900000 ;
    END
  END boot_addr_i[10]
  PIN boot_addr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.9865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 30.4197 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 162.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 48.6707 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 256.079 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 90.200000 0.000000 90.580000 0.900000 ;
    END
  END boot_addr_i[9]
  PIN boot_addr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5491 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 39.2037 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 209.552 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 73.0933 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 385.11 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 92.500000 0.000000 92.880000 0.900000 ;
    END
  END boot_addr_i[8]
  PIN boot_addr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9899 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.7885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.2776 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.088 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 94.2048 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 484.695 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 94.800000 0.000000 95.180000 0.900000 ;
    END
  END boot_addr_i[7]
  PIN boot_addr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.9569 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.6235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 56.5061 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 281.762 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 97.100000 0.000000 97.480000 0.900000 ;
    END
  END boot_addr_i[6]
  PIN boot_addr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7961 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.7015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.4134 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.0008 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 53.808 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 56.9434 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 298.053 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 99.400000 0.000000 99.780000 0.900000 ;
    END
  END boot_addr_i[5]
  PIN boot_addr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.5726 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.5258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 72.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 61.8473 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 327.168 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 101.700000 0.000000 102.080000 0.900000 ;
    END
  END boot_addr_i[4]
  PIN boot_addr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.0225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.151 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.824 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 73.0097 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 393.333 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 104.000000 0.000000 104.380000 0.900000 ;
    END
  END boot_addr_i[3]
  PIN boot_addr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4417 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.9295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.8912 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.968 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 30.0792 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 160.768 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 106.300000 0.000000 106.680000 0.900000 ;
    END
  END boot_addr_i[2]
  PIN boot_addr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3559 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.218 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.848 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 34.8848 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 190.032 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 108.600000 0.000000 108.980000 0.900000 ;
    END
  END boot_addr_i[1]
  PIN boot_addr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.2861 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.1515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.8088 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.784 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 58.3188 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 289.79 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 110.900000 0.000000 111.280000 0.900000 ;
    END
  END boot_addr_i[0]
  PIN instr_req_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4342 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.063 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 113.200000 0.000000 113.580000 0.900000 ;
    END
  END instr_req_o
  PIN instr_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.127 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.409 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 11.7306 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.8228 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.301829 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 115.500000 0.000000 115.880000 0.900000 ;
    END
  END instr_gnt_i
  PIN instr_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1054 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.183 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 10.2883 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.894 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 117.800000 0.000000 118.180000 0.900000 ;
    END
  END instr_rvalid_i
  PIN instr_addr_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7362 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 120.100000 0.000000 120.480000 0.900000 ;
    END
  END instr_addr_o[31]
  PIN instr_addr_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7664 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.596 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 122.400000 0.000000 122.780000 0.900000 ;
    END
  END instr_addr_o[30]
  PIN instr_addr_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.8872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.092 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 124.700000 0.000000 125.080000 0.900000 ;
    END
  END instr_addr_o[29]
  PIN instr_addr_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7954 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.751 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 127.000000 0.000000 127.380000 0.900000 ;
    END
  END instr_addr_o[28]
  PIN instr_addr_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.837 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.841 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 129.300000 0.000000 129.680000 0.900000 ;
    END
  END instr_addr_o[27]
  PIN instr_addr_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5949 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.2428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.432 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 131.600000 0.000000 131.980000 0.900000 ;
    END
  END instr_addr_o[26]
  PIN instr_addr_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5604 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 133.900000 0.000000 134.280000 0.900000 ;
    END
  END instr_addr_o[25]
  PIN instr_addr_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.9772 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.768 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 136.200000 0.000000 136.580000 0.900000 ;
    END
  END instr_addr_o[24]
  PIN instr_addr_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.7886 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 42.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 138.500000 0.000000 138.880000 0.900000 ;
    END
  END instr_addr_o[23]
  PIN instr_addr_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9366 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.457 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 140.800000 0.000000 141.180000 0.900000 ;
    END
  END instr_addr_o[22]
  PIN instr_addr_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0752 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.258 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 142.640000 0.000000 143.020000 0.900000 ;
    END
  END instr_addr_o[21]
  PIN instr_addr_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2274 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.675 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 144.940000 0.000000 145.320000 0.900000 ;
    END
  END instr_addr_o[20]
  PIN instr_addr_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4366 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.075 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 147.240000 0.000000 147.620000 0.900000 ;
    END
  END instr_addr_o[19]
  PIN instr_addr_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.623 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 149.540000 0.000000 149.920000 0.900000 ;
    END
  END instr_addr_o[18]
  PIN instr_addr_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.459 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 151.840000 0.000000 152.220000 0.900000 ;
    END
  END instr_addr_o[17]
  PIN instr_addr_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.5168 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 120.56 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 154.140000 0.000000 154.520000 0.900000 ;
    END
  END instr_addr_o[16]
  PIN instr_addr_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1203 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.6108 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99.728 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 156.440000 0.000000 156.820000 0.900000 ;
    END
  END instr_addr_o[15]
  PIN instr_addr_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6674 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.111 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 158.740000 0.000000 159.120000 0.900000 ;
    END
  END instr_addr_o[14]
  PIN instr_addr_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.875 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.149 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 161.040000 0.000000 161.420000 0.900000 ;
    END
  END instr_addr_o[13]
  PIN instr_addr_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.4336 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.92 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 163.340000 0.000000 163.720000 0.900000 ;
    END
  END instr_addr_o[12]
  PIN instr_addr_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5375 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.6878 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.472 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 165.640000 0.000000 166.020000 0.900000 ;
    END
  END instr_addr_o[11]
  PIN instr_addr_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.6765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.6378 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.872 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 167.940000 0.000000 168.320000 0.900000 ;
    END
  END instr_addr_o[10]
  PIN instr_addr_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.459 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 170.240000 0.000000 170.620000 0.900000 ;
    END
  END instr_addr_o[9]
  PIN instr_addr_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3822 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.685 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 172.540000 0.000000 172.920000 0.900000 ;
    END
  END instr_addr_o[8]
  PIN instr_addr_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3139 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.4808 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 174.840000 0.000000 175.220000 0.900000 ;
    END
  END instr_addr_o[7]
  PIN instr_addr_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3514 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.531 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 177.140000 0.000000 177.520000 0.900000 ;
    END
  END instr_addr_o[6]
  PIN instr_addr_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2347 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.0125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.6748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.736 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 179.440000 0.000000 179.820000 0.900000 ;
    END
  END instr_addr_o[5]
  PIN instr_addr_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.599 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 181.740000 0.000000 182.120000 0.900000 ;
    END
  END instr_addr_o[4]
  PIN instr_addr_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3233 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.1788 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.424 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 184.040000 0.000000 184.420000 0.900000 ;
    END
  END instr_addr_o[3]
  PIN instr_addr_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6034 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.791 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 186.340000 0.000000 186.720000 0.900000 ;
    END
  END instr_addr_o[2]
  PIN instr_addr_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1602 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.575 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 188.640000 0.000000 189.020000 0.900000 ;
    END
  END instr_addr_o[1]
  PIN instr_addr_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.755 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 190.940000 0.000000 191.320000 0.900000 ;
    END
  END instr_addr_o[0]
  PIN instr_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.168 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.6238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 78.464 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 93.8455 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 476.716 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.831217 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 193.240000 0.000000 193.620000 0.900000 ;
    END
  END instr_rdata_i[31]
  PIN instr_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7523 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.6005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.4038 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 66.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 73.2554 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 367.97 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.97672 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 195.540000 0.000000 195.920000 0.900000 ;
    END
  END instr_rdata_i[30]
  PIN instr_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7103 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.3905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.9268 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 60.8062 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 307.897 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.831217 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 197.840000 0.000000 198.220000 0.900000 ;
    END
  END instr_rdata_i[29]
  PIN instr_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3349 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.276 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.4648 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 77.616 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 87.9721 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 450.225 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32725 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 200.140000 0.000000 200.520000 0.900000 ;
    END
  END instr_rdata_i[28]
  PIN instr_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4507 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.9745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.9247 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.064 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met3  ;
    ANTENNAMAXAREACAR 45.304 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 220.486 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 202.440000 0.000000 202.820000 0.900000 ;
    END
  END instr_rdata_i[27]
  PIN instr_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.0225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.8386 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.08 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met3  ;
    ANTENNAMAXAREACAR 55.2591 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 272.981 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 204.740000 0.000000 205.120000 0.900000 ;
    END
  END instr_rdata_i[26]
  PIN instr_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9899 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.2356 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.7102 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 80.336 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 90.6075 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 477.243 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.36032 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 207.040000 0.000000 207.420000 0.900000 ;
    END
  END instr_rdata_i[25]
  PIN instr_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.9118 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.989 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met2  ;
    ANTENNAMAXAREACAR 39.9131 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 187.036 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.340000 0.000000 209.720000 0.900000 ;
    END
  END instr_rdata_i[24]
  PIN instr_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8213 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.5915 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 36.4873 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 169.05 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.4648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.616 LAYER met3  ;
    ANTENNAGATEAREA 0.378 LAYER met3  ;
    ANTENNAMAXAREACAR 43.0079 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 205.071 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 211.640000 0.000000 212.020000 0.900000 ;
    END
  END instr_rdata_i[23]
  PIN instr_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.2282 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.581 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met2  ;
    ANTENNAMAXAREACAR 22.6266 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 101.165 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 213.940000 0.000000 214.320000 0.900000 ;
    END
  END instr_rdata_i[22]
  PIN instr_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3559 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.9938 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.104 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met3  ;
    ANTENNAMAXAREACAR 50.3959 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 245.582 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.513757 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 216.240000 0.000000 216.620000 0.900000 ;
    END
  END instr_rdata_i[21]
  PIN instr_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.2166 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.621 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met2  ;
    ANTENNAMAXAREACAR 26.7739 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 121.304 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 218.540000 0.000000 218.920000 0.900000 ;
    END
  END instr_rdata_i[20]
  PIN instr_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.9786 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.559 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met2  ;
    ANTENNAMAXAREACAR 45.9115 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 216.795 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 220.840000 0.000000 221.220000 0.900000 ;
    END
  END instr_rdata_i[19]
  PIN instr_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.1026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.061 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met2  ;
    ANTENNAMAXAREACAR 28.8136 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 131.851 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 223.140000 0.000000 223.520000 0.900000 ;
    END
  END instr_rdata_i[18]
  PIN instr_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.3235 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.1025 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 36.0286 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 167.077 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.423 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.056 LAYER met3  ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 53.5802 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 262.538 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 55.3468 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 273.204 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 225.440000 0.000000 225.820000 0.900000 ;
    END
  END instr_rdata_i[17]
  PIN instr_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5444 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.335 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 31.3595 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 143.599 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.974603 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.757 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.504 LAYER met3  ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 46.2683 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 224.964 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.13333 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.0468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.72 LAYER met4  ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 54.3286 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 269.197 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.13333 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 227.740000 0.000000 228.120000 0.900000 ;
    END
  END instr_rdata_i[16]
  PIN instr_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.4974 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.163 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met2  ;
    ANTENNAMAXAREACAR 26.8015 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 122.128 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 230.040000 0.000000 230.420000 0.900000 ;
    END
  END instr_rdata_i[15]
  PIN instr_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2731 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.0965 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 30.8996 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 141.341 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 32.8909 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 155.69 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.1708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.048 LAYER met4  ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 54.5067 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 272.22 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 232.340000 0.000000 232.720000 0.900000 ;
    END
  END instr_rdata_i[14]
  PIN instr_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6426 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.879 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met2  ;
    ANTENNAMAXAREACAR 26.806 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 121.267 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 234.640000 0.000000 235.020000 0.900000 ;
    END
  END instr_rdata_i[13]
  PIN instr_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.0348 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met2  ;
    ANTENNAMAXAREACAR 28.2231 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 128.925 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 236.940000 0.000000 237.320000 0.900000 ;
    END
  END instr_rdata_i[12]
  PIN instr_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.265 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met2  ;
    ANTENNAMAXAREACAR 27.703 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 126.61 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.240000 0.000000 239.620000 0.900000 ;
    END
  END instr_rdata_i[11]
  PIN instr_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.4395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.5107 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.856 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met3  ;
    ANTENNAMAXAREACAR 28.9754 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 139.575 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 241.540000 0.000000 241.920000 0.900000 ;
    END
  END instr_rdata_i[10]
  PIN instr_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.0046 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.571 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met2  ;
    ANTENNAMAXAREACAR 33.5758 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 154.804 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 243.840000 0.000000 244.220000 0.900000 ;
    END
  END instr_rdata_i[9]
  PIN instr_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5949 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.229 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.6828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 52.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 50.8892 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 258.069 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.00979 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 246.140000 0.000000 246.520000 0.900000 ;
    END
  END instr_rdata_i[8]
  PIN instr_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3821 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.3547 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 109.024 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 75.3274 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 391.669 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 248.440000 0.000000 248.820000 0.900000 ;
    END
  END instr_rdata_i[7]
  PIN instr_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9417 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.5475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.4518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 50.88 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 49.9351 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 248.918 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.619577 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 250.740000 0.000000 251.120000 0.900000 ;
    END
  END instr_rdata_i[6]
  PIN instr_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0863 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.2705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.1708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 60.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 57.544 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 287.296 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.798148 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 253.040000 0.000000 253.420000 0.900000 ;
    END
  END instr_rdata_i[5]
  PIN instr_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1889 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.7796 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.432 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 103.23 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 536.501 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.67778 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 255.340000 0.000000 255.720000 0.900000 ;
    END
  END instr_rdata_i[4]
  PIN instr_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4847 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.5836 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 94.72 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 76.7382 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 390.5 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.798148 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 257.640000 0.000000 258.020000 0.900000 ;
    END
  END instr_rdata_i[3]
  PIN instr_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6497 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.197 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.7938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 68.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 64.621 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 324.099 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.798148 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 259.940000 0.000000 260.320000 0.900000 ;
    END
  END instr_rdata_i[2]
  PIN instr_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.351 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.788 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 95.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.0288 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 112.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 99.7382 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 512.048 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.619577 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 262.240000 0.000000 262.620000 0.900000 ;
    END
  END instr_rdata_i[1]
  PIN instr_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6989 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.1806 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 97.904 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 73.931 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 376.536 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.798148 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 264.540000 0.000000 264.920000 0.900000 ;
    END
  END instr_rdata_i[0]
  PIN data_req_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4342 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.063 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 266.840000 0.000000 267.220000 0.900000 ;
    END
  END data_req_o
  PIN data_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7899 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.5115 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 16.5739 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 79.4828 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.0696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.28 LAYER met3  ;
    ANTENNAGATEAREA 2.061 LAYER met3  ;
    ANTENNAMAXAREACAR 20.9745 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 103.394 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.550317 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.9618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.6 LAYER met4  ;
    ANTENNAGATEAREA 3.0555 LAYER met4  ;
    ANTENNAMAXAREACAR 22.2711 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 110.463 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.606888 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 269.140000 0.000000 269.520000 0.900000 ;
    END
  END data_gnt_i
  PIN data_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3092 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.933 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 17.0746 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 75.1438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.461484 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.586 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.592 LAYER met3  ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 25.8912 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 122.79 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.515032 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.4466 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.656 LAYER met4  ;
    ANTENNAGATEAREA 8.811 LAYER met4  ;
    ANTENNAMAXAREACAR 26.3959 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 125.589 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.515032 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 271.440000 0.000000 271.820000 0.900000 ;
    END
  END data_rvalid_i
  PIN data_we_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.6046 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.797 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 273.740000 0.000000 274.120000 0.900000 ;
    END
  END data_we_o
  PIN data_be_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4342 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.063 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 275.580000 0.000000 275.960000 0.900000 ;
    END
  END data_be_o[3]
  PIN data_be_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6034 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.791 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 277.880000 0.000000 278.260000 0.900000 ;
    END
  END data_be_o[2]
  PIN data_be_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.865 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.217 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 280.180000 0.000000 280.560000 0.900000 ;
    END
  END data_be_o[1]
  PIN data_be_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.651 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.029 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 282.480000 0.000000 282.860000 0.900000 ;
    END
  END data_be_o[0]
  PIN data_addr_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7829 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.7978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 127.392 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 284.780000 0.000000 285.160000 0.900000 ;
    END
  END data_addr_o[31]
  PIN data_addr_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6593 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.1355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.2008 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 124.208 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 287.080000 0.000000 287.460000 0.900000 ;
    END
  END data_addr_o[30]
  PIN data_addr_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9761 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.3948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.576 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 289.380000 0.000000 289.760000 0.900000 ;
    END
  END data_addr_o[29]
  PIN data_addr_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.9378 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 64.463 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 291.680000 0.000000 292.060000 0.900000 ;
    END
  END data_addr_o[28]
  PIN data_addr_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.5426 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.487 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 293.980000 0.000000 294.360000 0.900000 ;
    END
  END data_addr_o[27]
  PIN data_addr_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4885 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.2815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.1508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 102.608 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 296.280000 0.000000 296.660000 0.900000 ;
    END
  END data_addr_o[26]
  PIN data_addr_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.1945 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.8115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 298.580000 0.000000 298.960000 0.900000 ;
    END
  END data_addr_o[25]
  PIN data_addr_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8415 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.0465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.2448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 65.776 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 300.880000 0.000000 301.260000 0.900000 ;
    END
  END data_addr_o[24]
  PIN data_addr_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8931 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.0268 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 107.28 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 303.180000 0.000000 303.560000 0.900000 ;
    END
  END data_addr_o[23]
  PIN data_addr_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1245 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.5648 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 104.816 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 305.480000 0.000000 305.860000 0.900000 ;
    END
  END data_addr_o[22]
  PIN data_addr_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8473 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.0178 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 123.232 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 307.780000 0.000000 308.160000 0.900000 ;
    END
  END data_addr_o[21]
  PIN data_addr_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7829 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.2858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 135.328 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 310.080000 0.000000 310.460000 0.900000 ;
    END
  END data_addr_o[20]
  PIN data_addr_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2533 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.1055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.6628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 110.672 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 312.380000 0.000000 312.760000 0.900000 ;
    END
  END data_addr_o[19]
  PIN data_addr_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2609 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.1435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.8438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.304 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 314.680000 0.000000 315.060000 0.900000 ;
    END
  END data_addr_o[18]
  PIN data_addr_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6745 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.2115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.9418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 80.16 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 316.980000 0.000000 317.360000 0.900000 ;
    END
  END data_addr_o[17]
  PIN data_addr_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3525 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.6015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.3798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 66.496 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 319.280000 0.000000 319.660000 0.900000 ;
    END
  END data_addr_o[16]
  PIN data_addr_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2533 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.1055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.0068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 133.84 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 321.580000 0.000000 321.960000 0.900000 ;
    END
  END data_addr_o[15]
  PIN data_addr_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4818 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.301 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 323.880000 0.000000 324.260000 0.900000 ;
    END
  END data_addr_o[14]
  PIN data_addr_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6034 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.791 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 326.180000 0.000000 326.560000 0.900000 ;
    END
  END data_addr_o[13]
  PIN data_addr_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.651 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.029 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 328.480000 0.000000 328.860000 0.900000 ;
    END
  END data_addr_o[12]
  PIN data_addr_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4818 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.301 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 330.780000 0.000000 331.160000 0.900000 ;
    END
  END data_addr_o[11]
  PIN data_addr_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6442 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.113 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 333.080000 0.000000 333.460000 0.900000 ;
    END
  END data_addr_o[10]
  PIN data_addr_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9537 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.3708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.448 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 335.380000 0.000000 335.760000 0.900000 ;
    END
  END data_addr_o[9]
  PIN data_addr_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0467 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.0725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.8048 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 42.096 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 337.680000 0.000000 338.060000 0.900000 ;
    END
  END data_addr_o[8]
  PIN data_addr_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5491 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.1248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 81.136 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 339.980000 0.000000 340.360000 0.900000 ;
    END
  END data_addr_o[7]
  PIN data_addr_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5082 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.315 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 342.280000 0.000000 342.660000 0.900000 ;
    END
  END data_addr_o[6]
  PIN data_addr_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3807 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.056 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.0898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 107.616 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 344.580000 0.000000 344.960000 0.900000 ;
    END
  END data_addr_o[5]
  PIN data_addr_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.351 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 346.880000 0.000000 347.260000 0.900000 ;
    END
  END data_addr_o[4]
  PIN data_addr_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2991 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.3345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.5238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.264 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 349.180000 0.000000 349.560000 0.900000 ;
    END
  END data_addr_o[3]
  PIN data_addr_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.563 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.707 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 351.480000 0.000000 351.860000 0.900000 ;
    END
  END data_addr_o[2]
  PIN data_addr_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9746 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.765 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 353.780000 0.000000 354.160000 0.900000 ;
    END
  END data_addr_o[1]
  PIN data_addr_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.651 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.029 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 356.080000 0.000000 356.460000 0.900000 ;
    END
  END data_addr_o[0]
  PIN data_wdata_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.039 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.087 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 358.380000 0.000000 358.760000 0.900000 ;
    END
  END data_wdata_o[31]
  PIN data_wdata_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.431 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 360.680000 0.000000 361.060000 0.900000 ;
    END
  END data_wdata_o[30]
  PIN data_wdata_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.6266 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.025 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 362.980000 0.000000 363.360000 0.900000 ;
    END
  END data_wdata_o[29]
  PIN data_wdata_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4342 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.063 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 365.280000 0.000000 365.660000 0.900000 ;
    END
  END data_wdata_o[28]
  PIN data_wdata_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3349 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.2078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.912 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 367.580000 0.000000 367.960000 0.900000 ;
    END
  END data_wdata_o[27]
  PIN data_wdata_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.577 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 369.880000 0.000000 370.260000 0.900000 ;
    END
  END data_wdata_o[26]
  PIN data_wdata_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9606 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.695 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 372.180000 0.000000 372.560000 0.900000 ;
    END
  END data_wdata_o[25]
  PIN data_wdata_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.7988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.064 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 374.480000 0.000000 374.860000 0.900000 ;
    END
  END data_wdata_o[24]
  PIN data_wdata_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9746 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.765 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 376.780000 0.000000 377.160000 0.900000 ;
    END
  END data_wdata_o[23]
  PIN data_wdata_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.515 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.467 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 379.080000 0.000000 379.460000 0.900000 ;
    END
  END data_wdata_o[22]
  PIN data_wdata_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9102 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.443 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 381.380000 0.000000 381.760000 0.900000 ;
    END
  END data_wdata_o[21]
  PIN data_wdata_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.3882 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.833 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 383.680000 0.000000 384.060000 0.900000 ;
    END
  END data_wdata_o[20]
  PIN data_wdata_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4661 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.1695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.5368 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 385.980000 0.000000 386.360000 0.900000 ;
    END
  END data_wdata_o[19]
  PIN data_wdata_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6034 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.791 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 388.280000 0.000000 388.660000 0.900000 ;
    END
  END data_wdata_o[18]
  PIN data_wdata_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.039 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.087 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 390.580000 0.000000 390.960000 0.900000 ;
    END
  END data_wdata_o[17]
  PIN data_wdata_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5558 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.553 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 392.880000 0.000000 393.260000 0.900000 ;
    END
  END data_wdata_o[16]
  PIN data_wdata_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.039 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.087 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 395.180000 0.000000 395.560000 0.900000 ;
    END
  END data_wdata_o[15]
  PIN data_wdata_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.431 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 397.480000 0.000000 397.860000 0.900000 ;
    END
  END data_wdata_o[14]
  PIN data_wdata_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1338 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.561 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 399.780000 0.000000 400.160000 0.900000 ;
    END
  END data_wdata_o[13]
  PIN data_wdata_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.581 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.797 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 402.080000 0.000000 402.460000 0.900000 ;
    END
  END data_wdata_o[12]
  PIN data_wdata_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3807 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.2818 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 60.64 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 404.380000 0.000000 404.760000 0.900000 ;
    END
  END data_wdata_o[11]
  PIN data_wdata_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.7938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 68.704 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 406.680000 0.000000 407.060000 0.900000 ;
    END
  END data_wdata_o[10]
  PIN data_wdata_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.9512 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.638 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 408.520000 0.000000 408.900000 0.900000 ;
    END
  END data_wdata_o[9]
  PIN data_wdata_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7746 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.765 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 410.820000 0.000000 411.200000 0.900000 ;
    END
  END data_wdata_o[8]
  PIN data_wdata_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.039 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.087 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 413.120000 0.000000 413.500000 0.900000 ;
    END
  END data_wdata_o[7]
  PIN data_wdata_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6986 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.267 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 415.420000 0.000000 415.800000 0.900000 ;
    END
  END data_wdata_o[6]
  PIN data_wdata_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1678 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.731 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 417.720000 0.000000 418.100000 0.900000 ;
    END
  END data_wdata_o[5]
  PIN data_wdata_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1679 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.9488 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.864 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 420.020000 0.000000 420.400000 0.900000 ;
    END
  END data_wdata_o[4]
  PIN data_wdata_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6034 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.791 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 422.320000 0.000000 422.700000 0.900000 ;
    END
  END data_wdata_o[3]
  PIN data_wdata_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7798 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.673 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 424.620000 0.000000 425.000000 0.900000 ;
    END
  END data_wdata_o[2]
  PIN data_wdata_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1412 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.598 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 426.920000 0.000000 427.300000 0.900000 ;
    END
  END data_wdata_o[1]
  PIN data_wdata_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7966 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.757 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 429.220000 0.000000 429.600000 0.900000 ;
    END
  END data_wdata_o[0]
  PIN data_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4022 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.559 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 21.7027 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 90.1306 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 431.520000 0.000000 431.900000 0.900000 ;
    END
  END data_rdata_i[31]
  PIN data_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4618 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.965 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 22.5983 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 93.8963 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 433.820000 0.000000 434.200000 0.900000 ;
    END
  END data_rdata_i[30]
  PIN data_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.9494 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.305 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 22.6299 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 94.7798 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 436.120000 0.000000 436.500000 0.900000 ;
    END
  END data_rdata_i[29]
  PIN data_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4686 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.881 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 24.6519 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 104.006 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 438.420000 0.000000 438.800000 0.900000 ;
    END
  END data_rdata_i[28]
  PIN data_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9567 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.2785 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 24.8778 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 105.798 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.472349 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.621 LAYER met3  ;
    ANTENNAMAXAREACAR 25.2818 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 108.709 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.536761 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.9378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.472 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 34.5694 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 158.873 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 440.720000 0.000000 441.100000 0.900000 ;
    END
  END data_rdata_i[27]
  PIN data_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.5724 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.292 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 34.0573 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 150.889 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 443.020000 0.000000 443.400000 0.900000 ;
    END
  END data_rdata_i[26]
  PIN data_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4409 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.9155 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 9.9398 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.3869 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.230101 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met3  ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 29.5486 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 128.36 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 445.320000 0.000000 445.700000 0.900000 ;
    END
  END data_rdata_i[25]
  PIN data_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2272 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.631 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 6.93212 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 33.0212 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.1208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.448 LAYER met3  ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 30.4589 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 135.839 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 447.620000 0.000000 448.000000 0.900000 ;
    END
  END data_rdata_i[24]
  PIN data_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7498 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.297 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 22.2627 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 92.9304 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 449.920000 0.000000 450.300000 0.900000 ;
    END
  END data_rdata_i[23]
  PIN data_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.6906 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.129 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 16.1501 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 62.5389 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 452.220000 0.000000 452.600000 0.900000 ;
    END
  END data_rdata_i[22]
  PIN data_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.9278 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.305 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 19.3279 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.5576 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 454.520000 0.000000 454.900000 0.900000 ;
    END
  END data_rdata_i[21]
  PIN data_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8475 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.9685 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 6.16505 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.6626 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.171 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.712 LAYER met3  ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 14.5913 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 75.5455 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.7198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.976 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 30.6913 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 143.358 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 456.820000 0.000000 457.200000 0.900000 ;
    END
  END data_rdata_i[20]
  PIN data_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.6834 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.975 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 22.7849 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 95.5549 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 459.120000 0.000000 459.500000 0.900000 ;
    END
  END data_rdata_i[19]
  PIN data_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.6088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 30.384 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 30.8392 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 140.689 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.693603 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 461.420000 0.000000 461.800000 0.900000 ;
    END
  END data_rdata_i[18]
  PIN data_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.1286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.201 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 20.0475 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.8682 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 463.720000 0.000000 464.100000 0.900000 ;
    END
  END data_rdata_i[17]
  PIN data_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.831 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.703 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 31.4047 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 138.641 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 466.020000 0.000000 466.400000 0.900000 ;
    END
  END data_rdata_i[16]
  PIN data_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.43 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.58 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 17.1399 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 67.1587 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 468.320000 0.000000 468.700000 0.900000 ;
    END
  END data_rdata_i[15]
  PIN data_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.7735 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 6.53798 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.2889 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.826 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.872 LAYER met3  ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 14.2673 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 73.4545 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.7788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.624 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 46.144 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 226.466 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.884127 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 470.620000 0.000000 471.000000 0.900000 ;
    END
  END data_rdata_i[14]
  PIN data_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4105 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.54061 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.404 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 7.16081 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 36.3212 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.4596 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.392 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 47.3795 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 223.821 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 472.920000 0.000000 473.300000 0.900000 ;
    END
  END data_rdata_i[13]
  PIN data_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6387 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8065 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 8.56364 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.8364 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.091 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.952 LAYER met3  ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 14.8081 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 74.0828 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.7458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 68.448 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 46.9623 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 224.593 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 475.220000 0.000000 475.600000 0.900000 ;
    END
  END data_rdata_i[12]
  PIN data_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.8614 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.983 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 19.3454 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 78.5154 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 477.520000 0.000000 477.900000 0.900000 ;
    END
  END data_rdata_i[11]
  PIN data_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.052 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.873 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 8.82929 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 42.6091 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.568 LAYER met3  ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 20.2313 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 104.363 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.9488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.864 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 22.8401 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 118.906 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.636111 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 479.820000 0.000000 480.200000 0.900000 ;
    END
  END data_rdata_i[10]
  PIN data_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1674 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.503 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 19.5114 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 79.332 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 482.120000 0.000000 482.500000 0.900000 ;
    END
  END data_rdata_i[9]
  PIN data_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.7516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 47.616 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 20.7119 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 91.4806 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.515032 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 484.420000 0.000000 484.800000 0.900000 ;
    END
  END data_rdata_i[8]
  PIN data_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.4388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.144 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 49.3771 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 241.91 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.515032 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 486.720000 0.000000 487.100000 0.900000 ;
    END
  END data_rdata_i[7]
  PIN data_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.064 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.76 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 26.2611 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 112.778 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 489.020000 0.000000 489.400000 0.900000 ;
    END
  END data_rdata_i[6]
  PIN data_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9971 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.8245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.8784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 90.48 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 36.021 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 189.515 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.3408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 50.288 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 73.1032 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 362.249 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.38016 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 491.320000 0.000000 491.700000 0.900000 ;
    END
  END data_rdata_i[5]
  PIN data_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.0445 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.7075 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 32.797 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 144.521 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.65092 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.0048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.496 LAYER met3  ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 56.8998 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 273.699 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 493.620000 0.000000 494.000000 0.900000 ;
    END
  END data_rdata_i[4]
  PIN data_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.6853 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.8035 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 19.2527 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.4823 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.472349 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.6448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 94.576 LAYER met3  ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 42.8736 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 204.09 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 495.920000 0.000000 496.300000 0.900000 ;
    END
  END data_rdata_i[3]
  PIN data_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6803 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.0009 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.8 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met3  ;
    ANTENNAMAXAREACAR 30.9846 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 142.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.536761 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.3046 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 93.232 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 69.8551 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 349.904 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 498.220000 0.000000 498.600000 0.900000 ;
    END
  END data_rdata_i[2]
  PIN data_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.0166 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.641 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 17.0976 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 67.1185 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 500.520000 0.000000 500.900000 0.900000 ;
    END
  END data_rdata_i[1]
  PIN data_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9327 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.8864 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.856 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 6.5996 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 34.9253 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.8658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 53.088 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 31.4798 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 146.931 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 502.820000 0.000000 503.200000 0.900000 ;
    END
  END data_rdata_i[0]
  PIN data_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.120000 0.000000 505.500000 0.900000 ;
    END
  END data_err_i
  PIN irq_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2551 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.9965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.9671 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 1.7388 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.2116 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 255.088 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3643 LAYER met4  ;
    ANTENNAMAXAREACAR 47.2119 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 229.604 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.36411 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 507.420000 0.000000 507.800000 0.900000 ;
    END
  END irq_i
  PIN irq_id_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6602 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.193 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 21.3768 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 103.218 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 509.720000 0.000000 510.100000 0.900000 ;
    END
  END irq_id_i[4]
  PIN irq_id_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9438 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.611 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.10404 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 42.1273 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 512.020000 0.000000 512.400000 0.900000 ;
    END
  END irq_id_i[3]
  PIN irq_id_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5486 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.635 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 11.5477 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 54.3455 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 514.320000 0.000000 514.700000 0.900000 ;
    END
  END irq_id_i[2]
  PIN irq_id_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8794 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.289 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.84384 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.8263 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 516.620000 0.000000 517.000000 0.900000 ;
    END
  END irq_id_i[1]
  PIN irq_id_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8342 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.063 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 14.7246 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 69.9576 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 518.920000 0.000000 519.300000 0.900000 ;
    END
  END irq_id_i[0]
  PIN irq_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.1466 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.625 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 532.720000 0.000000 533.100000 0.900000 ;
    END
  END irq_ack_o
  PIN irq_id_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4818 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.301 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 521.220000 0.000000 521.600000 0.900000 ;
    END
  END irq_id_o[4]
  PIN irq_id_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9102 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.443 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 523.520000 0.000000 523.900000 0.900000 ;
    END
  END irq_id_o[3]
  PIN irq_id_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6106 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.945 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 525.820000 0.000000 526.200000 0.900000 ;
    END
  END irq_id_o[2]
  PIN irq_id_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.563 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.707 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 528.120000 0.000000 528.500000 0.900000 ;
    END
  END irq_id_o[1]
  PIN irq_id_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9102 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.443 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 530.420000 0.000000 530.800000 0.900000 ;
    END
  END irq_id_o[0]
  PIN debug_req_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4599 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.737 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 39.1758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 211.76 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 92.7283 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 489.766 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.36032 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 535.020000 0.000000 535.400000 0.900000 ;
    END
  END debug_req_i
  PIN fetch_enable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.6293 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.6215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.7412 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.168 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 37.1065 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 195.119 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 537.320000 0.000000 537.700000 0.900000 ;
    END
  END fetch_enable_i
  PIN ext_perf_counters_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.3305 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.4915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 56.1592 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 301.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9936 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.24 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 74.9385 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 387.448 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 539.160000 0.000000 539.540000 0.900000 ;
    END
  END ext_perf_counters_i
  PIN eFPGA_operand_a_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 9.840000 550.160000 10.220000 ;
    END
  END eFPGA_operand_a_o[31]
  PIN eFPGA_operand_a_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 58.0668 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 310.16 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 12.890000 550.160000 13.270000 ;
    END
  END eFPGA_operand_a_o[30]
  PIN eFPGA_operand_a_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.0906 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.0374 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 150.944 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 15.940000 550.160000 16.320000 ;
    END
  END eFPGA_operand_a_o[29]
  PIN eFPGA_operand_a_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5546 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.7356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 164.864 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 18.990000 550.160000 19.370000 ;
    END
  END eFPGA_operand_a_o[28]
  PIN eFPGA_operand_a_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4526 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.8622 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 134.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 22.040000 550.160000 22.420000 ;
    END
  END eFPGA_operand_a_o[27]
  PIN eFPGA_operand_a_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 45.5784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 243.08 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 25.090000 550.160000 25.470000 ;
    END
  END eFPGA_operand_a_o[26]
  PIN eFPGA_operand_a_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1256 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.2618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 119.2 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 28.750000 550.160000 29.130000 ;
    END
  END eFPGA_operand_a_o[25]
  PIN eFPGA_operand_a_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 47.8734 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 255.32 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 31.800000 550.160000 32.180000 ;
    END
  END eFPGA_operand_a_o[24]
  PIN eFPGA_operand_a_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2326 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.1956 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 97.984 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 34.850000 550.160000 35.230000 ;
    END
  END eFPGA_operand_a_o[23]
  PIN eFPGA_operand_a_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 31.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 169.208 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 37.900000 550.160000 38.280000 ;
    END
  END eFPGA_operand_a_o[22]
  PIN eFPGA_operand_a_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 47.3184 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 252.36 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 40.950000 550.160000 41.330000 ;
    END
  END eFPGA_operand_a_o[21]
  PIN eFPGA_operand_a_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 39.1374 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 208.728 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 44.000000 550.160000 44.380000 ;
    END
  END eFPGA_operand_a_o[20]
  PIN eFPGA_operand_a_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.5256 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.9248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.736 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 47.050000 550.160000 47.430000 ;
    END
  END eFPGA_operand_a_o[19]
  PIN eFPGA_operand_a_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.8672 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.424 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 50.710000 550.160000 51.090000 ;
    END
  END eFPGA_operand_a_o[18]
  PIN eFPGA_operand_a_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.7146 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.752 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 53.760000 550.160000 54.140000 ;
    END
  END eFPGA_operand_a_o[17]
  PIN eFPGA_operand_a_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 38.8024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 207.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.6808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.768 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 56.810000 550.160000 57.190000 ;
    END
  END eFPGA_operand_a_o[16]
  PIN eFPGA_operand_a_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.1436 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.1436 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 71.04 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 59.860000 550.160000 60.240000 ;
    END
  END eFPGA_operand_a_o[15]
  PIN eFPGA_operand_a_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 37.9264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 202.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.3612 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 131.808 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 62.910000 550.160000 63.290000 ;
    END
  END eFPGA_operand_a_o[14]
  PIN eFPGA_operand_a_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.1766 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 235.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.7796 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.432 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 66.570000 550.160000 66.950000 ;
    END
  END eFPGA_operand_a_o[13]
  PIN eFPGA_operand_a_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.4736 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 173.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.3408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 50.288 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 69.620000 550.160000 70.000000 ;
    END
  END eFPGA_operand_a_o[12]
  PIN eFPGA_operand_a_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 70.7394 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 377.272 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 72.670000 550.160000 73.050000 ;
    END
  END eFPGA_operand_a_o[11]
  PIN eFPGA_operand_a_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 57.2992 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 306.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 75.720000 550.160000 76.100000 ;
    END
  END eFPGA_operand_a_o[10]
  PIN eFPGA_operand_a_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.2096 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 155.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.4084 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 62.256 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 78.770000 550.160000 79.150000 ;
    END
  END eFPGA_operand_a_o[9]
  PIN eFPGA_operand_a_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 60.9162 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 325.352 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 81.820000 550.160000 82.200000 ;
    END
  END eFPGA_operand_a_o[8]
  PIN eFPGA_operand_a_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 85.480000 550.160000 85.860000 ;
    END
  END eFPGA_operand_a_o[7]
  PIN eFPGA_operand_a_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2776 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.6296 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.632 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 88.530000 550.160000 88.910000 ;
    END
  END eFPGA_operand_a_o[6]
  PIN eFPGA_operand_a_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 91.580000 550.160000 91.960000 ;
    END
  END eFPGA_operand_a_o[5]
  PIN eFPGA_operand_a_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4846 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.936 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 94.630000 550.160000 95.010000 ;
    END
  END eFPGA_operand_a_o[4]
  PIN eFPGA_operand_a_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 79.0554 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 421.624 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 97.680000 550.160000 98.060000 ;
    END
  END eFPGA_operand_a_o[3]
  PIN eFPGA_operand_a_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.6096 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 120.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.1066 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.176 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 100.730000 550.160000 101.110000 ;
    END
  END eFPGA_operand_a_o[2]
  PIN eFPGA_operand_a_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.852 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 106.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.2876 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.808 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 104.390000 550.160000 104.770000 ;
    END
  END eFPGA_operand_a_o[1]
  PIN eFPGA_operand_a_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 64.9066 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 346.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 107.440000 550.160000 107.820000 ;
    END
  END eFPGA_operand_a_o[0]
  PIN eFPGA_operand_b_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.0552 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 160.76 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 110.490000 550.160000 110.870000 ;
    END
  END eFPGA_operand_b_o[31]
  PIN eFPGA_operand_b_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.1304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.024 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 113.540000 550.160000 113.920000 ;
    END
  END eFPGA_operand_b_o[30]
  PIN eFPGA_operand_b_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.2416 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 129.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 116.590000 550.160000 116.970000 ;
    END
  END eFPGA_operand_b_o[29]
  PIN eFPGA_operand_b_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.9776 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 111.872 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 119.640000 550.160000 120.020000 ;
    END
  END eFPGA_operand_b_o[28]
  PIN eFPGA_operand_b_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.2064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.096 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 122.690000 550.160000 123.070000 ;
    END
  END eFPGA_operand_b_o[27]
  PIN eFPGA_operand_b_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 23.1774 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.608 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 126.350000 550.160000 126.730000 ;
    END
  END eFPGA_operand_b_o[26]
  PIN eFPGA_operand_b_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 129.400000 550.160000 129.780000 ;
    END
  END eFPGA_operand_b_o[25]
  PIN eFPGA_operand_b_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.8714 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.976 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 132.450000 550.160000 132.830000 ;
    END
  END eFPGA_operand_b_o[24]
  PIN eFPGA_operand_b_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.3784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.68 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 135.500000 550.160000 135.880000 ;
    END
  END eFPGA_operand_b_o[23]
  PIN eFPGA_operand_b_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 138.550000 550.160000 138.930000 ;
    END
  END eFPGA_operand_b_o[22]
  PIN eFPGA_operand_b_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 141.600000 550.160000 141.980000 ;
    END
  END eFPGA_operand_b_o[21]
  PIN eFPGA_operand_b_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 145.260000 550.160000 145.640000 ;
    END
  END eFPGA_operand_b_o[20]
  PIN eFPGA_operand_b_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 28.9254 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 154.264 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 148.310000 550.160000 148.690000 ;
    END
  END eFPGA_operand_b_o[19]
  PIN eFPGA_operand_b_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 28.5084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 152.04 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 151.360000 550.160000 151.740000 ;
    END
  END eFPGA_operand_b_o[18]
  PIN eFPGA_operand_b_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 154.410000 550.160000 154.790000 ;
    END
  END eFPGA_operand_b_o[17]
  PIN eFPGA_operand_b_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 157.460000 550.160000 157.840000 ;
    END
  END eFPGA_operand_b_o[16]
  PIN eFPGA_operand_b_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 160.510000 550.160000 160.890000 ;
    END
  END eFPGA_operand_b_o[15]
  PIN eFPGA_operand_b_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.7334 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 164.170000 550.160000 164.550000 ;
    END
  END eFPGA_operand_b_o[14]
  PIN eFPGA_operand_b_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 167.220000 550.160000 167.600000 ;
    END
  END eFPGA_operand_b_o[13]
  PIN eFPGA_operand_b_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 170.270000 550.160000 170.650000 ;
    END
  END eFPGA_operand_b_o[12]
  PIN eFPGA_operand_b_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 45.2994 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 241.592 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 173.320000 550.160000 173.700000 ;
    END
  END eFPGA_operand_b_o[11]
  PIN eFPGA_operand_b_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.5666 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.0736 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 92 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 176.370000 550.160000 176.750000 ;
    END
  END eFPGA_operand_b_o[10]
  PIN eFPGA_operand_b_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.3476 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 184.128 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 179.420000 550.160000 179.800000 ;
    END
  END eFPGA_operand_b_o[9]
  PIN eFPGA_operand_b_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 44.1504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 235.464 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 183.080000 550.160000 183.460000 ;
    END
  END eFPGA_operand_b_o[8]
  PIN eFPGA_operand_b_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 37.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 201.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 186.130000 550.160000 186.510000 ;
    END
  END eFPGA_operand_b_o[7]
  PIN eFPGA_operand_b_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 42.5712 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 227.512 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 189.180000 550.160000 189.560000 ;
    END
  END eFPGA_operand_b_o[6]
  PIN eFPGA_operand_b_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4846 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.1928 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.832 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 192.230000 550.160000 192.610000 ;
    END
  END eFPGA_operand_b_o[5]
  PIN eFPGA_operand_b_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 195.280000 550.160000 195.660000 ;
    END
  END eFPGA_operand_b_o[4]
  PIN eFPGA_operand_b_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 40.4326 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 215.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.6808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.768 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 198.940000 550.160000 199.320000 ;
    END
  END eFPGA_operand_b_o[3]
  PIN eFPGA_operand_b_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4406 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.4978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.792 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 201.990000 550.160000 202.370000 ;
    END
  END eFPGA_operand_b_o[2]
  PIN eFPGA_operand_b_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 41.3424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 220.488 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 205.040000 550.160000 205.420000 ;
    END
  END eFPGA_operand_b_o[1]
  PIN eFPGA_operand_b_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 41.3364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 220.456 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 208.090000 550.160000 208.470000 ;
    END
  END eFPGA_operand_b_o[0]
  PIN eFPGA_result_a_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4774 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 69.1547 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 343.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 211.140000 550.160000 211.520000 ;
    END
  END eFPGA_result_a_i[31]
  PIN eFPGA_result_a_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.288 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 65.6873 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 324.994 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 214.190000 550.160000 214.570000 ;
    END
  END eFPGA_result_a_i[30]
  PIN eFPGA_result_a_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8944 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.432 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 72.7572 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 361.895 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 217.850000 550.160000 218.230000 ;
    END
  END eFPGA_result_a_i[29]
  PIN eFPGA_result_a_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.864 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 14.5899 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 68.4929 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 220.900000 550.160000 221.280000 ;
    END
  END eFPGA_result_a_i[28]
  PIN eFPGA_result_a_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 19.8141 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 93.499 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 223.950000 550.160000 224.330000 ;
    END
  END eFPGA_result_a_i[27]
  PIN eFPGA_result_a_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 20.0743 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 94.1253 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 227.000000 550.160000 227.380000 ;
    END
  END eFPGA_result_a_i[26]
  PIN eFPGA_result_a_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.064 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 62.0905 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 309.984 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 230.050000 550.160000 230.430000 ;
    END
  END eFPGA_result_a_i[25]
  PIN eFPGA_result_a_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 63.0368 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 309.414 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 233.100000 550.160000 233.480000 ;
    END
  END eFPGA_result_a_i[24]
  PIN eFPGA_result_a_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 63.1224 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 310.376 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 236.760000 550.160000 237.140000 ;
    END
  END eFPGA_result_a_i[23]
  PIN eFPGA_result_a_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.392 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 12.6986 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 58.9253 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 239.810000 550.160000 240.190000 ;
    END
  END eFPGA_result_a_i[22]
  PIN eFPGA_result_a_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0184 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.9378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.472 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 35.5523 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 186.505 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 242.860000 550.160000 243.240000 ;
    END
  END eFPGA_result_a_i[21]
  PIN eFPGA_result_a_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.92 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 12.122 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 55.4101 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 245.910000 550.160000 246.290000 ;
    END
  END eFPGA_result_a_i[20]
  PIN eFPGA_result_a_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4846 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.8418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 68.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 63.4707 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 333.18 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 248.960000 550.160000 249.340000 ;
    END
  END eFPGA_result_a_i[19]
  PIN eFPGA_result_a_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.4188 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 98.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 77.9224 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 412.145 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 252.010000 550.160000 252.390000 ;
    END
  END eFPGA_result_a_i[18]
  PIN eFPGA_result_a_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.224 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 64.059 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 317.846 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 255.670000 550.160000 256.050000 ;
    END
  END eFPGA_result_a_i[17]
  PIN eFPGA_result_a_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.864 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 22.0234 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 105.77 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 258.720000 550.160000 259.100000 ;
    END
  END eFPGA_result_a_i[16]
  PIN eFPGA_result_a_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 10.9366 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 49.5475 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 261.770000 550.160000 262.150000 ;
    END
  END eFPGA_result_a_i[15]
  PIN eFPGA_result_a_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.736 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 16.779 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 81.5758 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 264.820000 550.160000 265.200000 ;
    END
  END eFPGA_result_a_i[14]
  PIN eFPGA_result_a_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.92 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 12.2109 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 56.004 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 267.870000 550.160000 268.250000 ;
    END
  END eFPGA_result_a_i[13]
  PIN eFPGA_result_a_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.864 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 13.6154 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 63.7697 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 270.920000 550.160000 271.300000 ;
    END
  END eFPGA_result_a_i[12]
  PIN eFPGA_result_a_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6864 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.656 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 11.9782 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 54.9899 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 274.580000 550.160000 274.960000 ;
    END
  END eFPGA_result_a_i[11]
  PIN eFPGA_result_a_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6864 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.656 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 11.697 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 53.802 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 277.630000 550.160000 278.010000 ;
    END
  END eFPGA_result_a_i[10]
  PIN eFPGA_result_a_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.584 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 22.8719 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 113.77 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 280.680000 550.160000 281.060000 ;
    END
  END eFPGA_result_a_i[9]
  PIN eFPGA_result_a_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.92 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 12.4711 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 57.305 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 283.730000 550.160000 284.110000 ;
    END
  END eFPGA_result_a_i[8]
  PIN eFPGA_result_a_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0184 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.76 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 16.6061 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 79.9596 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 286.780000 550.160000 287.160000 ;
    END
  END eFPGA_result_a_i[7]
  PIN eFPGA_result_a_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.92 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 13.6364 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 63.1313 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 289.830000 550.160000 290.210000 ;
    END
  END eFPGA_result_a_i[6]
  PIN eFPGA_result_a_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.584 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 19.857 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 98.6949 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 293.490000 550.160000 293.870000 ;
    END
  END eFPGA_result_a_i[5]
  PIN eFPGA_result_a_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6184 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.96 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 49.8246 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 246.861 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 296.540000 550.160000 296.920000 ;
    END
  END eFPGA_result_a_i[4]
  PIN eFPGA_result_a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2044 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.752 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 51.1895 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 253.127 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 299.590000 550.160000 299.970000 ;
    END
  END eFPGA_result_a_i[3]
  PIN eFPGA_result_a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.7796 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.432 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 69.9782 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 370.525 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 302.640000 550.160000 303.020000 ;
    END
  END eFPGA_result_a_i[2]
  PIN eFPGA_result_a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.288 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 47.9313 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 236.214 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 305.690000 550.160000 306.070000 ;
    END
  END eFPGA_result_a_i[1]
  PIN eFPGA_result_a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.5888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 88.944 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 77.0044 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 405.648 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 308.740000 550.160000 309.120000 ;
    END
  END eFPGA_result_a_i[0]
  PIN eFPGA_result_b_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.264 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 57.1349 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 278.54 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 312.400000 550.160000 312.780000 ;
    END
  END eFPGA_result_b_i[31]
  PIN eFPGA_result_b_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.424 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 62.2032 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 305.944 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 315.450000 550.160000 315.830000 ;
    END
  END eFPGA_result_b_i[30]
  PIN eFPGA_result_b_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.6764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.936 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 74.3667 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 372.968 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 318.500000 550.160000 318.880000 ;
    END
  END eFPGA_result_b_i[29]
  PIN eFPGA_result_b_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.376 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 47.4286 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 227.087 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 321.550000 550.160000 321.930000 ;
    END
  END eFPGA_result_b_i[28]
  PIN eFPGA_result_b_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5614 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.656 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 63.681 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 313.944 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 324.600000 550.160000 324.980000 ;
    END
  END eFPGA_result_b_i[27]
  PIN eFPGA_result_b_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9054 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.824 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 63.2159 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 307.238 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 327.650000 550.160000 328.030000 ;
    END
  END eFPGA_result_b_i[26]
  PIN eFPGA_result_b_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0654 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.344 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 80.8476 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 401.111 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 331.310000 550.160000 331.690000 ;
    END
  END eFPGA_result_b_i[25]
  PIN eFPGA_result_b_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 60.3603 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 296.127 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 334.360000 550.160000 334.740000 ;
    END
  END eFPGA_result_b_i[24]
  PIN eFPGA_result_b_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.624 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 67.1873 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 332.452 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 337.410000 550.160000 337.790000 ;
    END
  END eFPGA_result_b_i[23]
  PIN eFPGA_result_b_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.304 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 71.7413 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 357.048 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 340.460000 550.160000 340.840000 ;
    END
  END eFPGA_result_b_i[22]
  PIN eFPGA_result_b_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6544 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.152 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 67.2635 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 332.103 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 343.510000 550.160000 343.890000 ;
    END
  END eFPGA_result_b_i[21]
  PIN eFPGA_result_b_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5954 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 59.681 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 291.389 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 346.560000 550.160000 346.940000 ;
    END
  END eFPGA_result_b_i[20]
  PIN eFPGA_result_b_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8294 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.752 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 58.7159 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 287.183 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 350.220000 550.160000 350.600000 ;
    END
  END eFPGA_result_b_i[19]
  PIN eFPGA_result_b_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 57.1968 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 279.214 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 353.270000 550.160000 353.650000 ;
    END
  END eFPGA_result_b_i[18]
  PIN eFPGA_result_b_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.9414 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 80.6151 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 402.802 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 356.320000 550.160000 356.700000 ;
    END
  END eFPGA_result_b_i[17]
  PIN eFPGA_result_b_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 65.4611 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 323.262 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 359.370000 550.160000 359.750000 ;
    END
  END eFPGA_result_b_i[16]
  PIN eFPGA_result_b_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6544 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.152 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 67.0746 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 331.159 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 362.420000 550.160000 362.800000 ;
    END
  END eFPGA_result_b_i[15]
  PIN eFPGA_result_b_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 28.4381 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 121.524 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 365.470000 550.160000 365.850000 ;
    END
  END eFPGA_result_b_i[14]
  PIN eFPGA_result_b_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9624 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.128 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 96.5762 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 463.444 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 369.130000 550.160000 369.510000 ;
    END
  END eFPGA_result_b_i[13]
  PIN eFPGA_result_b_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3826 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.4978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.792 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 79.0921 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 417.627 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 372.180000 550.160000 372.560000 ;
    END
  END eFPGA_result_b_i[12]
  PIN eFPGA_result_b_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.5598 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.392 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 88.6476 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 451.683 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 375.230000 550.160000 375.610000 ;
    END
  END eFPGA_result_b_i[11]
  PIN eFPGA_result_b_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6524 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 48.0794 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 223.429 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 378.280000 550.160000 378.660000 ;
    END
  END eFPGA_result_b_i[10]
  PIN eFPGA_result_b_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 100.51 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 480.349 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 381.330000 550.160000 381.710000 ;
    END
  END eFPGA_result_b_i[9]
  PIN eFPGA_result_b_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 55.9429 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 257.516 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 384.380000 550.160000 384.760000 ;
    END
  END eFPGA_result_b_i[8]
  PIN eFPGA_result_b_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.914 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.144 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 80.9857 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 414.159 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 388.040000 550.160000 388.420000 ;
    END
  END eFPGA_result_b_i[7]
  PIN eFPGA_result_b_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.3222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.984 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.3168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 50.16 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 112.429 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 584.214 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 391.090000 550.160000 391.470000 ;
    END
  END eFPGA_result_b_i[6]
  PIN eFPGA_result_b_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6524 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 36.8159 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 169.484 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 394.140000 550.160000 394.520000 ;
    END
  END eFPGA_result_b_i[5]
  PIN eFPGA_result_b_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 95.2825 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 470.738 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 397.190000 550.160000 397.570000 ;
    END
  END eFPGA_result_b_i[4]
  PIN eFPGA_result_b_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8374 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.128 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 97.4976 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 484.294 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 400.240000 550.160000 400.620000 ;
    END
  END eFPGA_result_b_i[3]
  PIN eFPGA_result_b_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 71.0159 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 339.183 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 403.290000 550.160000 403.670000 ;
    END
  END eFPGA_result_b_i[2]
  PIN eFPGA_result_b_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6174 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.288 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 111.44 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 555.532 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 406.340000 550.160000 406.720000 ;
    END
  END eFPGA_result_b_i[1]
  PIN eFPGA_result_b_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.784 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 111.8 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 557.579 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 410.000000 550.160000 410.380000 ;
    END
  END eFPGA_result_b_i[0]
  PIN eFPGA_result_c_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.0138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 64.544 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 100.435 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 520.279 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 413.050000 550.160000 413.430000 ;
    END
  END eFPGA_result_c_i[31]
  PIN eFPGA_result_c_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.904 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 80.9263 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 406.667 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 416.100000 550.160000 416.480000 ;
    END
  END eFPGA_result_c_i[30]
  PIN eFPGA_result_c_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.4648 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 61.616 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 97.184 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 503.749 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 419.150000 550.160000 419.530000 ;
    END
  END eFPGA_result_c_i[29]
  PIN eFPGA_result_c_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 16.4261 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 80.1131 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 422.200000 550.160000 422.580000 ;
    END
  END eFPGA_result_c_i[28]
  PIN eFPGA_result_c_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.0106 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.664 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 67.7449 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 364.687 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 425.250000 550.160000 425.630000 ;
    END
  END eFPGA_result_c_i[27]
  PIN eFPGA_result_c_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.864 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 26.8883 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 132.941 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 428.910000 550.160000 429.290000 ;
    END
  END eFPGA_result_c_i[26]
  PIN eFPGA_result_c_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0664 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 90.5844 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 453.471 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 431.960000 550.160000 432.340000 ;
    END
  END eFPGA_result_c_i[25]
  PIN eFPGA_result_c_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 17.5913 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 85.9394 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 435.010000 550.160000 435.390000 ;
    END
  END eFPGA_result_c_i[24]
  PIN eFPGA_result_c_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0664 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 15.4584 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 78.0727 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 438.060000 550.160000 438.440000 ;
    END
  END eFPGA_result_c_i[23]
  PIN eFPGA_result_c_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0832 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 22.8313 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 120.941 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 441.110000 550.160000 441.490000 ;
    END
  END eFPGA_result_c_i[22]
  PIN eFPGA_result_c_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9624 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.128 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 15.5339 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 76.7394 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 444.160000 550.160000 444.540000 ;
    END
  END eFPGA_result_c_i[21]
  PIN eFPGA_result_c_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.912 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 82.0414 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 411.992 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 447.820000 550.160000 448.200000 ;
    END
  END eFPGA_result_c_i[20]
  PIN eFPGA_result_c_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.1598 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 53.5178 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 280.699 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 450.870000 550.160000 451.250000 ;
    END
  END eFPGA_result_c_i[19]
  PIN eFPGA_result_c_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 70.1473 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 348.521 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 453.920000 550.160000 454.300000 ;
    END
  END eFPGA_result_c_i[18]
  PIN eFPGA_result_c_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4846 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.7568 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 73.84 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 60.3497 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 322.174 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 456.970000 550.160000 457.350000 ;
    END
  END eFPGA_result_c_i[17]
  PIN eFPGA_result_c_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.92 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 82.8051 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 412.529 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 460.020000 550.160000 460.400000 ;
    END
  END eFPGA_result_c_i[16]
  PIN eFPGA_result_c_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6524 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 23.0887 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 115.394 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 463.070000 550.160000 463.450000 ;
    END
  END eFPGA_result_c_i[15]
  PIN eFPGA_result_c_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.89395 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.0268 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.28 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 84.5901 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 444.962 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 466.730000 550.160000 467.110000 ;
    END
  END eFPGA_result_c_i[14]
  PIN eFPGA_result_c_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.2326 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.0948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.976 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 34.6919 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 184.028 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 469.780000 550.160000 470.160000 ;
    END
  END eFPGA_result_c_i[13]
  PIN eFPGA_result_c_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5694 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.0378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 80.672 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 77.9121 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 412.238 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 472.830000 550.160000 473.210000 ;
    END
  END eFPGA_result_c_i[12]
  PIN eFPGA_result_c_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 18.2927 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 88.7717 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 475.880000 550.160000 476.260000 ;
    END
  END eFPGA_result_c_i[11]
  PIN eFPGA_result_c_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.28 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 87.8644 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 438.194 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 478.930000 550.160000 479.310000 ;
    END
  END eFPGA_result_c_i[10]
  PIN eFPGA_result_c_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.7924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 81.3909 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 437.709 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 481.980000 550.160000 482.360000 ;
    END
  END eFPGA_result_c_i[9]
  PIN eFPGA_result_c_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.92 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 52.7566 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 260.707 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 485.640000 550.160000 486.020000 ;
    END
  END eFPGA_result_c_i[8]
  PIN eFPGA_result_c_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.864 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 13.883 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 68.5131 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 488.690000 550.160000 489.070000 ;
    END
  END eFPGA_result_c_i[7]
  PIN eFPGA_result_c_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.92 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 12.1566 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 59.6162 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 491.740000 550.160000 492.120000 ;
    END
  END eFPGA_result_c_i[6]
  PIN eFPGA_result_c_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9624 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.128 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 13.2362 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 65.596 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 494.790000 550.160000 495.170000 ;
    END
  END eFPGA_result_c_i[5]
  PIN eFPGA_result_c_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 14.2863 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 71.8343 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 497.840000 550.160000 498.220000 ;
    END
  END eFPGA_result_c_i[4]
  PIN eFPGA_result_c_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.488 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 95.0935 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 476.388 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 500.890000 550.160000 501.270000 ;
    END
  END eFPGA_result_c_i[3]
  PIN eFPGA_result_c_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.32 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 93.7343 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 468.792 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 504.550000 550.160000 504.930000 ;
    END
  END eFPGA_result_c_i[2]
  PIN eFPGA_result_c_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5154 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 15.9558 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 83.7495 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 507.600000 550.160000 507.980000 ;
    END
  END eFPGA_result_c_i[1]
  PIN eFPGA_result_c_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 12.0176 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 57.7131 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 510.650000 550.160000 511.030000 ;
    END
  END eFPGA_result_c_i[0]
  PIN eFPGA_write_strobe_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.3784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.68 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 513.700000 550.160000 514.080000 ;
    END
  END eFPGA_write_strobe_o
  PIN eFPGA_fpga_done_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.584 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met3  ;
    ANTENNAMAXAREACAR 19.1224 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 79.4493 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.472349 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 516.750000 550.160000 517.130000 ;
    END
  END eFPGA_fpga_done_i
  PIN eFPGA_en_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.0664 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.016 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 519.800000 550.160000 520.180000 ;
    END
  END eFPGA_en_o
  PIN eFPGA_operator_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 523.460000 550.160000 523.840000 ;
    END
  END eFPGA_operator_o[1]
  PIN eFPGA_operator_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 526.510000 550.160000 526.890000 ;
    END
  END eFPGA_operator_o[0]
  PIN eFPGA_delay_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 529.560000 550.160000 529.940000 ;
    END
  END eFPGA_delay_o[3]
  PIN eFPGA_delay_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.3764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.336 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 532.610000 550.160000 532.990000 ;
    END
  END eFPGA_delay_o[2]
  PIN eFPGA_delay_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 535.660000 550.160000 536.040000 ;
    END
  END eFPGA_delay_o[1]
  PIN eFPGA_delay_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.2044 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.752 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 538.710000 550.160000 539.090000 ;
    END
  END eFPGA_delay_o[0]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 548.960000 541.960000 550.160000 543.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 541.960000 1.200000 543.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 548.960000 5.430000 550.160000 6.630000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 5.430000 1.200000 6.630000 ;
    END
    PORT
      LAYER met4 ;
        RECT 543.400000 548.580000 544.600000 549.780000 ;
    END
    PORT
      LAYER met4 ;
        RECT 543.400000 0.000000 544.600000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 5.560000 548.580000 6.760000 549.780000 ;
    END
    PORT
      LAYER met4 ;
        RECT 5.560000 0.000000 6.760000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 5.430000 550.160000 6.630000 ;
        RECT 0.000000 541.960000 550.160000 543.160000 ;
        RECT 5.560000 9.620000 6.760000 10.100000 ;
        RECT 5.560000 15.060000 6.760000 15.540000 ;
        RECT 12.120000 9.620000 13.320000 10.100000 ;
        RECT 12.120000 15.060000 13.320000 15.540000 ;
        RECT 5.560000 20.500000 6.760000 20.980000 ;
        RECT 12.120000 20.500000 13.320000 20.980000 ;
        RECT 5.560000 25.940000 6.760000 26.420000 ;
        RECT 5.560000 31.380000 6.760000 31.860000 ;
        RECT 12.120000 31.380000 13.320000 31.860000 ;
        RECT 12.120000 25.940000 13.320000 26.420000 ;
        RECT 57.120000 31.380000 58.320000 31.860000 ;
        RECT 57.120000 25.940000 58.320000 26.420000 ;
        RECT 57.120000 20.500000 58.320000 20.980000 ;
        RECT 57.120000 15.060000 58.320000 15.540000 ;
        RECT 57.120000 9.620000 58.320000 10.100000 ;
        RECT 5.560000 36.820000 6.760000 37.300000 ;
        RECT 5.560000 42.260000 6.760000 42.740000 ;
        RECT 12.120000 42.260000 13.320000 42.740000 ;
        RECT 12.120000 36.820000 13.320000 37.300000 ;
        RECT 5.560000 47.700000 6.760000 48.180000 ;
        RECT 12.120000 47.700000 13.320000 48.180000 ;
        RECT 5.560000 53.140000 6.760000 53.620000 ;
        RECT 5.560000 58.580000 6.760000 59.060000 ;
        RECT 12.120000 58.580000 13.320000 59.060000 ;
        RECT 12.120000 53.140000 13.320000 53.620000 ;
        RECT 5.560000 64.020000 6.760000 64.500000 ;
        RECT 12.120000 64.020000 13.320000 64.500000 ;
        RECT 57.120000 47.700000 58.320000 48.180000 ;
        RECT 57.120000 42.260000 58.320000 42.740000 ;
        RECT 57.120000 36.820000 58.320000 37.300000 ;
        RECT 57.120000 58.580000 58.320000 59.060000 ;
        RECT 57.120000 53.140000 58.320000 53.620000 ;
        RECT 57.120000 64.020000 58.320000 64.500000 ;
        RECT 102.120000 9.620000 103.320000 10.100000 ;
        RECT 102.120000 15.060000 103.320000 15.540000 ;
        RECT 102.120000 20.500000 103.320000 20.980000 ;
        RECT 102.120000 25.940000 103.320000 26.420000 ;
        RECT 102.120000 31.380000 103.320000 31.860000 ;
        RECT 102.120000 64.020000 103.320000 64.500000 ;
        RECT 102.120000 36.820000 103.320000 37.300000 ;
        RECT 102.120000 42.260000 103.320000 42.740000 ;
        RECT 102.120000 47.700000 103.320000 48.180000 ;
        RECT 102.120000 53.140000 103.320000 53.620000 ;
        RECT 102.120000 58.580000 103.320000 59.060000 ;
        RECT 5.560000 69.460000 6.760000 69.940000 ;
        RECT 5.560000 74.900000 6.760000 75.380000 ;
        RECT 12.120000 74.900000 13.320000 75.380000 ;
        RECT 12.120000 69.460000 13.320000 69.940000 ;
        RECT 5.560000 80.340000 6.760000 80.820000 ;
        RECT 12.120000 80.340000 13.320000 80.820000 ;
        RECT 5.560000 85.780000 6.760000 86.260000 ;
        RECT 12.120000 85.780000 13.320000 86.260000 ;
        RECT 12.120000 91.220000 13.320000 91.700000 ;
        RECT 5.560000 91.220000 6.760000 91.700000 ;
        RECT 5.560000 96.660000 6.760000 97.140000 ;
        RECT 5.560000 102.100000 6.760000 102.580000 ;
        RECT 12.120000 96.660000 13.320000 97.140000 ;
        RECT 12.120000 102.100000 13.320000 102.580000 ;
        RECT 57.120000 80.340000 58.320000 80.820000 ;
        RECT 57.120000 74.900000 58.320000 75.380000 ;
        RECT 57.120000 69.460000 58.320000 69.940000 ;
        RECT 57.120000 85.780000 58.320000 86.260000 ;
        RECT 57.120000 91.220000 58.320000 91.700000 ;
        RECT 57.120000 96.660000 58.320000 97.140000 ;
        RECT 57.120000 102.100000 58.320000 102.580000 ;
        RECT 5.560000 107.540000 6.760000 108.020000 ;
        RECT 12.120000 107.540000 13.320000 108.020000 ;
        RECT 5.560000 112.980000 6.760000 113.460000 ;
        RECT 5.560000 118.420000 6.760000 118.900000 ;
        RECT 12.120000 118.420000 13.320000 118.900000 ;
        RECT 12.120000 112.980000 13.320000 113.460000 ;
        RECT 5.560000 123.860000 6.760000 124.340000 ;
        RECT 12.120000 123.860000 13.320000 124.340000 ;
        RECT 5.560000 129.300000 6.760000 129.780000 ;
        RECT 5.560000 134.740000 6.760000 135.220000 ;
        RECT 12.120000 129.300000 13.320000 129.780000 ;
        RECT 12.120000 134.740000 13.320000 135.220000 ;
        RECT 57.120000 118.420000 58.320000 118.900000 ;
        RECT 57.120000 112.980000 58.320000 113.460000 ;
        RECT 57.120000 107.540000 58.320000 108.020000 ;
        RECT 57.120000 129.300000 58.320000 129.780000 ;
        RECT 57.120000 123.860000 58.320000 124.340000 ;
        RECT 57.120000 134.740000 58.320000 135.220000 ;
        RECT 102.120000 80.340000 103.320000 80.820000 ;
        RECT 102.120000 74.900000 103.320000 75.380000 ;
        RECT 102.120000 69.460000 103.320000 69.940000 ;
        RECT 102.120000 85.780000 103.320000 86.260000 ;
        RECT 102.120000 91.220000 103.320000 91.700000 ;
        RECT 102.120000 96.660000 103.320000 97.140000 ;
        RECT 102.120000 102.100000 103.320000 102.580000 ;
        RECT 102.120000 134.740000 103.320000 135.220000 ;
        RECT 102.120000 129.300000 103.320000 129.780000 ;
        RECT 102.120000 123.860000 103.320000 124.340000 ;
        RECT 102.120000 107.540000 103.320000 108.020000 ;
        RECT 102.120000 112.980000 103.320000 113.460000 ;
        RECT 102.120000 118.420000 103.320000 118.900000 ;
        RECT 147.120000 31.380000 148.320000 31.860000 ;
        RECT 147.120000 25.940000 148.320000 26.420000 ;
        RECT 147.120000 20.500000 148.320000 20.980000 ;
        RECT 147.120000 15.060000 148.320000 15.540000 ;
        RECT 147.120000 9.620000 148.320000 10.100000 ;
        RECT 192.120000 31.380000 193.320000 31.860000 ;
        RECT 192.120000 25.940000 193.320000 26.420000 ;
        RECT 192.120000 15.060000 193.320000 15.540000 ;
        RECT 192.120000 9.620000 193.320000 10.100000 ;
        RECT 192.120000 20.500000 193.320000 20.980000 ;
        RECT 147.120000 47.700000 148.320000 48.180000 ;
        RECT 147.120000 42.260000 148.320000 42.740000 ;
        RECT 147.120000 36.820000 148.320000 37.300000 ;
        RECT 147.120000 58.580000 148.320000 59.060000 ;
        RECT 147.120000 53.140000 148.320000 53.620000 ;
        RECT 147.120000 64.020000 148.320000 64.500000 ;
        RECT 192.120000 47.700000 193.320000 48.180000 ;
        RECT 192.120000 42.260000 193.320000 42.740000 ;
        RECT 192.120000 36.820000 193.320000 37.300000 ;
        RECT 192.120000 58.580000 193.320000 59.060000 ;
        RECT 192.120000 53.140000 193.320000 53.620000 ;
        RECT 192.120000 64.020000 193.320000 64.500000 ;
        RECT 237.120000 9.620000 238.320000 10.100000 ;
        RECT 237.120000 15.060000 238.320000 15.540000 ;
        RECT 237.120000 20.500000 238.320000 20.980000 ;
        RECT 237.120000 25.940000 238.320000 26.420000 ;
        RECT 237.120000 31.380000 238.320000 31.860000 ;
        RECT 237.120000 36.820000 238.320000 37.300000 ;
        RECT 237.120000 42.260000 238.320000 42.740000 ;
        RECT 237.120000 47.700000 238.320000 48.180000 ;
        RECT 237.120000 64.020000 238.320000 64.500000 ;
        RECT 237.120000 53.140000 238.320000 53.620000 ;
        RECT 237.120000 58.580000 238.320000 59.060000 ;
        RECT 147.120000 80.340000 148.320000 80.820000 ;
        RECT 147.120000 74.900000 148.320000 75.380000 ;
        RECT 147.120000 69.460000 148.320000 69.940000 ;
        RECT 147.120000 96.660000 148.320000 97.140000 ;
        RECT 147.120000 85.780000 148.320000 86.260000 ;
        RECT 147.120000 91.220000 148.320000 91.700000 ;
        RECT 147.120000 102.100000 148.320000 102.580000 ;
        RECT 192.120000 80.340000 193.320000 80.820000 ;
        RECT 192.120000 74.900000 193.320000 75.380000 ;
        RECT 192.120000 69.460000 193.320000 69.940000 ;
        RECT 192.120000 85.780000 193.320000 86.260000 ;
        RECT 192.120000 91.220000 193.320000 91.700000 ;
        RECT 192.120000 96.660000 193.320000 97.140000 ;
        RECT 192.120000 102.100000 193.320000 102.580000 ;
        RECT 147.120000 118.420000 148.320000 118.900000 ;
        RECT 147.120000 112.980000 148.320000 113.460000 ;
        RECT 147.120000 107.540000 148.320000 108.020000 ;
        RECT 147.120000 129.300000 148.320000 129.780000 ;
        RECT 147.120000 123.860000 148.320000 124.340000 ;
        RECT 147.120000 134.740000 148.320000 135.220000 ;
        RECT 192.120000 118.420000 193.320000 118.900000 ;
        RECT 192.120000 112.980000 193.320000 113.460000 ;
        RECT 192.120000 107.540000 193.320000 108.020000 ;
        RECT 192.120000 129.300000 193.320000 129.780000 ;
        RECT 192.120000 123.860000 193.320000 124.340000 ;
        RECT 192.120000 134.740000 193.320000 135.220000 ;
        RECT 237.120000 80.340000 238.320000 80.820000 ;
        RECT 237.120000 74.900000 238.320000 75.380000 ;
        RECT 237.120000 69.460000 238.320000 69.940000 ;
        RECT 237.120000 85.780000 238.320000 86.260000 ;
        RECT 237.120000 91.220000 238.320000 91.700000 ;
        RECT 237.120000 96.660000 238.320000 97.140000 ;
        RECT 237.120000 102.100000 238.320000 102.580000 ;
        RECT 237.120000 107.540000 238.320000 108.020000 ;
        RECT 237.120000 112.980000 238.320000 113.460000 ;
        RECT 237.120000 118.420000 238.320000 118.900000 ;
        RECT 237.120000 134.740000 238.320000 135.220000 ;
        RECT 237.120000 129.300000 238.320000 129.780000 ;
        RECT 237.120000 123.860000 238.320000 124.340000 ;
        RECT 12.120000 145.620000 13.320000 146.100000 ;
        RECT 5.560000 145.620000 6.760000 146.100000 ;
        RECT 12.120000 140.180000 13.320000 140.660000 ;
        RECT 5.560000 140.180000 6.760000 140.660000 ;
        RECT 5.560000 151.060000 6.760000 151.540000 ;
        RECT 12.120000 151.060000 13.320000 151.540000 ;
        RECT 5.560000 156.500000 6.760000 156.980000 ;
        RECT 5.560000 161.940000 6.760000 162.420000 ;
        RECT 12.120000 156.500000 13.320000 156.980000 ;
        RECT 12.120000 161.940000 13.320000 162.420000 ;
        RECT 5.560000 167.380000 6.760000 167.860000 ;
        RECT 12.120000 167.380000 13.320000 167.860000 ;
        RECT 57.120000 145.620000 58.320000 146.100000 ;
        RECT 57.120000 140.180000 58.320000 140.660000 ;
        RECT 57.120000 151.060000 58.320000 151.540000 ;
        RECT 57.120000 156.500000 58.320000 156.980000 ;
        RECT 57.120000 161.940000 58.320000 162.420000 ;
        RECT 57.120000 167.380000 58.320000 167.860000 ;
        RECT 5.560000 172.820000 6.760000 173.300000 ;
        RECT 5.560000 178.260000 6.760000 178.740000 ;
        RECT 12.120000 178.260000 13.320000 178.740000 ;
        RECT 12.120000 172.820000 13.320000 173.300000 ;
        RECT 5.560000 183.700000 6.760000 184.180000 ;
        RECT 12.120000 183.700000 13.320000 184.180000 ;
        RECT 5.560000 189.140000 6.760000 189.620000 ;
        RECT 12.120000 194.580000 13.320000 195.060000 ;
        RECT 12.120000 189.140000 13.320000 189.620000 ;
        RECT 5.560000 194.580000 6.760000 195.060000 ;
        RECT 5.560000 200.020000 6.760000 200.500000 ;
        RECT 5.560000 205.460000 6.760000 205.940000 ;
        RECT 12.120000 200.020000 13.320000 200.500000 ;
        RECT 12.120000 205.460000 13.320000 205.940000 ;
        RECT 57.120000 183.700000 58.320000 184.180000 ;
        RECT 57.120000 178.260000 58.320000 178.740000 ;
        RECT 57.120000 172.820000 58.320000 173.300000 ;
        RECT 57.120000 194.580000 58.320000 195.060000 ;
        RECT 57.120000 189.140000 58.320000 189.620000 ;
        RECT 57.120000 200.020000 58.320000 200.500000 ;
        RECT 57.120000 205.460000 58.320000 205.940000 ;
        RECT 102.120000 145.620000 103.320000 146.100000 ;
        RECT 102.120000 140.180000 103.320000 140.660000 ;
        RECT 102.120000 151.060000 103.320000 151.540000 ;
        RECT 102.120000 156.500000 103.320000 156.980000 ;
        RECT 102.120000 161.940000 103.320000 162.420000 ;
        RECT 102.120000 167.380000 103.320000 167.860000 ;
        RECT 102.120000 205.460000 103.320000 205.940000 ;
        RECT 102.120000 200.020000 103.320000 200.500000 ;
        RECT 102.120000 194.580000 103.320000 195.060000 ;
        RECT 102.120000 172.820000 103.320000 173.300000 ;
        RECT 102.120000 178.260000 103.320000 178.740000 ;
        RECT 102.120000 183.700000 103.320000 184.180000 ;
        RECT 102.120000 189.140000 103.320000 189.620000 ;
        RECT 5.560000 210.900000 6.760000 211.380000 ;
        RECT 12.120000 210.900000 13.320000 211.380000 ;
        RECT 5.560000 216.340000 6.760000 216.820000 ;
        RECT 5.560000 221.780000 6.760000 222.260000 ;
        RECT 12.120000 221.780000 13.320000 222.260000 ;
        RECT 12.120000 216.340000 13.320000 216.820000 ;
        RECT 5.560000 227.220000 6.760000 227.700000 ;
        RECT 12.120000 227.220000 13.320000 227.700000 ;
        RECT 5.560000 232.660000 6.760000 233.140000 ;
        RECT 5.560000 238.100000 6.760000 238.580000 ;
        RECT 12.120000 238.100000 13.320000 238.580000 ;
        RECT 12.120000 232.660000 13.320000 233.140000 ;
        RECT 57.120000 221.780000 58.320000 222.260000 ;
        RECT 57.120000 216.340000 58.320000 216.820000 ;
        RECT 57.120000 210.900000 58.320000 211.380000 ;
        RECT 57.120000 227.220000 58.320000 227.700000 ;
        RECT 57.120000 232.660000 58.320000 233.140000 ;
        RECT 57.120000 238.100000 58.320000 238.580000 ;
        RECT 12.120000 248.980000 13.320000 249.460000 ;
        RECT 5.560000 248.980000 6.760000 249.460000 ;
        RECT 12.120000 243.540000 13.320000 244.020000 ;
        RECT 5.560000 243.540000 6.760000 244.020000 ;
        RECT 5.560000 254.420000 6.760000 254.900000 ;
        RECT 12.120000 254.420000 13.320000 254.900000 ;
        RECT 5.560000 259.860000 6.760000 260.340000 ;
        RECT 5.560000 265.300000 6.760000 265.780000 ;
        RECT 12.120000 265.300000 13.320000 265.780000 ;
        RECT 12.120000 259.860000 13.320000 260.340000 ;
        RECT 5.560000 270.740000 6.760000 271.220000 ;
        RECT 12.120000 270.740000 13.320000 271.220000 ;
        RECT 57.120000 254.420000 58.320000 254.900000 ;
        RECT 57.120000 248.980000 58.320000 249.460000 ;
        RECT 57.120000 243.540000 58.320000 244.020000 ;
        RECT 57.120000 265.300000 58.320000 265.780000 ;
        RECT 57.120000 259.860000 58.320000 260.340000 ;
        RECT 57.120000 270.740000 58.320000 271.220000 ;
        RECT 102.120000 221.780000 103.320000 222.260000 ;
        RECT 102.120000 216.340000 103.320000 216.820000 ;
        RECT 102.120000 210.900000 103.320000 211.380000 ;
        RECT 102.120000 227.220000 103.320000 227.700000 ;
        RECT 102.120000 232.660000 103.320000 233.140000 ;
        RECT 102.120000 238.100000 103.320000 238.580000 ;
        RECT 102.120000 270.740000 103.320000 271.220000 ;
        RECT 102.120000 265.300000 103.320000 265.780000 ;
        RECT 102.120000 243.540000 103.320000 244.020000 ;
        RECT 102.120000 248.980000 103.320000 249.460000 ;
        RECT 102.120000 254.420000 103.320000 254.900000 ;
        RECT 102.120000 259.860000 103.320000 260.340000 ;
        RECT 147.120000 140.180000 148.320000 140.660000 ;
        RECT 147.120000 145.620000 148.320000 146.100000 ;
        RECT 147.120000 151.060000 148.320000 151.540000 ;
        RECT 147.120000 167.380000 148.320000 167.860000 ;
        RECT 147.120000 156.500000 148.320000 156.980000 ;
        RECT 147.120000 161.940000 148.320000 162.420000 ;
        RECT 192.120000 140.180000 193.320000 140.660000 ;
        RECT 192.120000 145.620000 193.320000 146.100000 ;
        RECT 192.120000 151.060000 193.320000 151.540000 ;
        RECT 192.120000 156.500000 193.320000 156.980000 ;
        RECT 192.120000 161.940000 193.320000 162.420000 ;
        RECT 192.120000 167.380000 193.320000 167.860000 ;
        RECT 147.120000 183.700000 148.320000 184.180000 ;
        RECT 147.120000 178.260000 148.320000 178.740000 ;
        RECT 147.120000 172.820000 148.320000 173.300000 ;
        RECT 147.120000 194.580000 148.320000 195.060000 ;
        RECT 147.120000 189.140000 148.320000 189.620000 ;
        RECT 147.120000 200.020000 148.320000 200.500000 ;
        RECT 147.120000 205.460000 148.320000 205.940000 ;
        RECT 192.120000 183.700000 193.320000 184.180000 ;
        RECT 192.120000 178.260000 193.320000 178.740000 ;
        RECT 192.120000 172.820000 193.320000 173.300000 ;
        RECT 192.120000 194.580000 193.320000 195.060000 ;
        RECT 192.120000 189.140000 193.320000 189.620000 ;
        RECT 192.120000 200.020000 193.320000 200.500000 ;
        RECT 192.120000 205.460000 193.320000 205.940000 ;
        RECT 237.120000 145.620000 238.320000 146.100000 ;
        RECT 237.120000 140.180000 238.320000 140.660000 ;
        RECT 237.120000 151.060000 238.320000 151.540000 ;
        RECT 237.120000 156.500000 238.320000 156.980000 ;
        RECT 237.120000 161.940000 238.320000 162.420000 ;
        RECT 237.120000 167.380000 238.320000 167.860000 ;
        RECT 237.120000 172.820000 238.320000 173.300000 ;
        RECT 237.120000 178.260000 238.320000 178.740000 ;
        RECT 237.120000 183.700000 238.320000 184.180000 ;
        RECT 237.120000 205.460000 238.320000 205.940000 ;
        RECT 237.120000 200.020000 238.320000 200.500000 ;
        RECT 237.120000 194.580000 238.320000 195.060000 ;
        RECT 237.120000 189.140000 238.320000 189.620000 ;
        RECT 147.120000 221.780000 148.320000 222.260000 ;
        RECT 147.120000 216.340000 148.320000 216.820000 ;
        RECT 147.120000 210.900000 148.320000 211.380000 ;
        RECT 147.120000 238.100000 148.320000 238.580000 ;
        RECT 147.120000 227.220000 148.320000 227.700000 ;
        RECT 147.120000 232.660000 148.320000 233.140000 ;
        RECT 192.120000 221.780000 193.320000 222.260000 ;
        RECT 192.120000 216.340000 193.320000 216.820000 ;
        RECT 192.120000 210.900000 193.320000 211.380000 ;
        RECT 192.120000 227.220000 193.320000 227.700000 ;
        RECT 192.120000 232.660000 193.320000 233.140000 ;
        RECT 192.120000 238.100000 193.320000 238.580000 ;
        RECT 147.120000 254.420000 148.320000 254.900000 ;
        RECT 147.120000 248.980000 148.320000 249.460000 ;
        RECT 147.120000 243.540000 148.320000 244.020000 ;
        RECT 147.120000 265.300000 148.320000 265.780000 ;
        RECT 147.120000 259.860000 148.320000 260.340000 ;
        RECT 147.120000 270.740000 148.320000 271.220000 ;
        RECT 192.120000 254.420000 193.320000 254.900000 ;
        RECT 192.120000 248.980000 193.320000 249.460000 ;
        RECT 192.120000 243.540000 193.320000 244.020000 ;
        RECT 192.120000 265.300000 193.320000 265.780000 ;
        RECT 192.120000 259.860000 193.320000 260.340000 ;
        RECT 192.120000 270.740000 193.320000 271.220000 ;
        RECT 237.120000 221.780000 238.320000 222.260000 ;
        RECT 237.120000 216.340000 238.320000 216.820000 ;
        RECT 237.120000 210.900000 238.320000 211.380000 ;
        RECT 237.120000 227.220000 238.320000 227.700000 ;
        RECT 237.120000 232.660000 238.320000 233.140000 ;
        RECT 237.120000 238.100000 238.320000 238.580000 ;
        RECT 237.120000 243.540000 238.320000 244.020000 ;
        RECT 237.120000 248.980000 238.320000 249.460000 ;
        RECT 237.120000 254.420000 238.320000 254.900000 ;
        RECT 237.120000 270.740000 238.320000 271.220000 ;
        RECT 237.120000 265.300000 238.320000 265.780000 ;
        RECT 237.120000 259.860000 238.320000 260.340000 ;
        RECT 282.120000 31.380000 283.320000 31.860000 ;
        RECT 282.120000 25.940000 283.320000 26.420000 ;
        RECT 282.120000 20.500000 283.320000 20.980000 ;
        RECT 282.120000 15.060000 283.320000 15.540000 ;
        RECT 282.120000 9.620000 283.320000 10.100000 ;
        RECT 327.120000 31.380000 328.320000 31.860000 ;
        RECT 327.120000 25.940000 328.320000 26.420000 ;
        RECT 327.120000 20.500000 328.320000 20.980000 ;
        RECT 327.120000 15.060000 328.320000 15.540000 ;
        RECT 327.120000 9.620000 328.320000 10.100000 ;
        RECT 282.120000 47.700000 283.320000 48.180000 ;
        RECT 282.120000 42.260000 283.320000 42.740000 ;
        RECT 282.120000 36.820000 283.320000 37.300000 ;
        RECT 282.120000 58.580000 283.320000 59.060000 ;
        RECT 282.120000 53.140000 283.320000 53.620000 ;
        RECT 282.120000 64.020000 283.320000 64.500000 ;
        RECT 327.120000 47.700000 328.320000 48.180000 ;
        RECT 327.120000 42.260000 328.320000 42.740000 ;
        RECT 327.120000 36.820000 328.320000 37.300000 ;
        RECT 327.120000 58.580000 328.320000 59.060000 ;
        RECT 327.120000 53.140000 328.320000 53.620000 ;
        RECT 327.120000 64.020000 328.320000 64.500000 ;
        RECT 372.120000 20.500000 373.320000 20.980000 ;
        RECT 372.120000 9.620000 373.320000 10.100000 ;
        RECT 372.120000 15.060000 373.320000 15.540000 ;
        RECT 372.120000 25.940000 373.320000 26.420000 ;
        RECT 372.120000 31.380000 373.320000 31.860000 ;
        RECT 372.120000 36.820000 373.320000 37.300000 ;
        RECT 372.120000 42.260000 373.320000 42.740000 ;
        RECT 372.120000 47.700000 373.320000 48.180000 ;
        RECT 372.120000 64.020000 373.320000 64.500000 ;
        RECT 372.120000 53.140000 373.320000 53.620000 ;
        RECT 372.120000 58.580000 373.320000 59.060000 ;
        RECT 282.120000 80.340000 283.320000 80.820000 ;
        RECT 282.120000 74.900000 283.320000 75.380000 ;
        RECT 282.120000 69.460000 283.320000 69.940000 ;
        RECT 282.120000 96.660000 283.320000 97.140000 ;
        RECT 282.120000 85.780000 283.320000 86.260000 ;
        RECT 282.120000 91.220000 283.320000 91.700000 ;
        RECT 282.120000 102.100000 283.320000 102.580000 ;
        RECT 327.120000 80.340000 328.320000 80.820000 ;
        RECT 327.120000 74.900000 328.320000 75.380000 ;
        RECT 327.120000 69.460000 328.320000 69.940000 ;
        RECT 327.120000 85.780000 328.320000 86.260000 ;
        RECT 327.120000 91.220000 328.320000 91.700000 ;
        RECT 327.120000 96.660000 328.320000 97.140000 ;
        RECT 327.120000 102.100000 328.320000 102.580000 ;
        RECT 282.120000 118.420000 283.320000 118.900000 ;
        RECT 282.120000 112.980000 283.320000 113.460000 ;
        RECT 282.120000 107.540000 283.320000 108.020000 ;
        RECT 282.120000 129.300000 283.320000 129.780000 ;
        RECT 282.120000 123.860000 283.320000 124.340000 ;
        RECT 282.120000 134.740000 283.320000 135.220000 ;
        RECT 327.120000 118.420000 328.320000 118.900000 ;
        RECT 327.120000 112.980000 328.320000 113.460000 ;
        RECT 327.120000 107.540000 328.320000 108.020000 ;
        RECT 327.120000 129.300000 328.320000 129.780000 ;
        RECT 327.120000 123.860000 328.320000 124.340000 ;
        RECT 327.120000 134.740000 328.320000 135.220000 ;
        RECT 372.120000 80.340000 373.320000 80.820000 ;
        RECT 372.120000 74.900000 373.320000 75.380000 ;
        RECT 372.120000 69.460000 373.320000 69.940000 ;
        RECT 372.120000 85.780000 373.320000 86.260000 ;
        RECT 372.120000 91.220000 373.320000 91.700000 ;
        RECT 372.120000 96.660000 373.320000 97.140000 ;
        RECT 372.120000 102.100000 373.320000 102.580000 ;
        RECT 372.120000 107.540000 373.320000 108.020000 ;
        RECT 372.120000 112.980000 373.320000 113.460000 ;
        RECT 372.120000 118.420000 373.320000 118.900000 ;
        RECT 372.120000 134.740000 373.320000 135.220000 ;
        RECT 372.120000 129.300000 373.320000 129.780000 ;
        RECT 372.120000 123.860000 373.320000 124.340000 ;
        RECT 417.120000 31.380000 418.320000 31.860000 ;
        RECT 417.120000 25.940000 418.320000 26.420000 ;
        RECT 417.120000 20.500000 418.320000 20.980000 ;
        RECT 417.120000 15.060000 418.320000 15.540000 ;
        RECT 417.120000 9.620000 418.320000 10.100000 ;
        RECT 462.120000 31.380000 463.320000 31.860000 ;
        RECT 462.120000 25.940000 463.320000 26.420000 ;
        RECT 462.120000 20.500000 463.320000 20.980000 ;
        RECT 462.120000 15.060000 463.320000 15.540000 ;
        RECT 462.120000 9.620000 463.320000 10.100000 ;
        RECT 417.120000 47.700000 418.320000 48.180000 ;
        RECT 417.120000 42.260000 418.320000 42.740000 ;
        RECT 417.120000 36.820000 418.320000 37.300000 ;
        RECT 417.120000 58.580000 418.320000 59.060000 ;
        RECT 417.120000 53.140000 418.320000 53.620000 ;
        RECT 417.120000 64.020000 418.320000 64.500000 ;
        RECT 462.120000 47.700000 463.320000 48.180000 ;
        RECT 462.120000 42.260000 463.320000 42.740000 ;
        RECT 462.120000 36.820000 463.320000 37.300000 ;
        RECT 462.120000 58.580000 463.320000 59.060000 ;
        RECT 462.120000 53.140000 463.320000 53.620000 ;
        RECT 462.120000 64.020000 463.320000 64.500000 ;
        RECT 507.120000 31.380000 508.320000 31.860000 ;
        RECT 507.120000 25.940000 508.320000 26.420000 ;
        RECT 507.120000 20.500000 508.320000 20.980000 ;
        RECT 507.120000 15.060000 508.320000 15.540000 ;
        RECT 507.120000 9.620000 508.320000 10.100000 ;
        RECT 543.400000 15.060000 544.600000 15.540000 ;
        RECT 543.400000 9.620000 544.600000 10.100000 ;
        RECT 543.400000 31.380000 544.600000 31.860000 ;
        RECT 543.400000 25.940000 544.600000 26.420000 ;
        RECT 543.400000 20.500000 544.600000 20.980000 ;
        RECT 507.120000 36.820000 508.320000 37.300000 ;
        RECT 507.120000 42.260000 508.320000 42.740000 ;
        RECT 507.120000 47.700000 508.320000 48.180000 ;
        RECT 507.120000 64.020000 508.320000 64.500000 ;
        RECT 507.120000 58.580000 508.320000 59.060000 ;
        RECT 507.120000 53.140000 508.320000 53.620000 ;
        RECT 543.400000 47.700000 544.600000 48.180000 ;
        RECT 543.400000 42.260000 544.600000 42.740000 ;
        RECT 543.400000 36.820000 544.600000 37.300000 ;
        RECT 543.400000 64.020000 544.600000 64.500000 ;
        RECT 543.400000 58.580000 544.600000 59.060000 ;
        RECT 543.400000 53.140000 544.600000 53.620000 ;
        RECT 417.120000 80.340000 418.320000 80.820000 ;
        RECT 417.120000 74.900000 418.320000 75.380000 ;
        RECT 417.120000 69.460000 418.320000 69.940000 ;
        RECT 417.120000 96.660000 418.320000 97.140000 ;
        RECT 417.120000 85.780000 418.320000 86.260000 ;
        RECT 417.120000 91.220000 418.320000 91.700000 ;
        RECT 417.120000 102.100000 418.320000 102.580000 ;
        RECT 462.120000 80.340000 463.320000 80.820000 ;
        RECT 462.120000 74.900000 463.320000 75.380000 ;
        RECT 462.120000 69.460000 463.320000 69.940000 ;
        RECT 462.120000 85.780000 463.320000 86.260000 ;
        RECT 462.120000 91.220000 463.320000 91.700000 ;
        RECT 462.120000 96.660000 463.320000 97.140000 ;
        RECT 462.120000 102.100000 463.320000 102.580000 ;
        RECT 417.120000 118.420000 418.320000 118.900000 ;
        RECT 417.120000 112.980000 418.320000 113.460000 ;
        RECT 417.120000 107.540000 418.320000 108.020000 ;
        RECT 417.120000 129.300000 418.320000 129.780000 ;
        RECT 417.120000 123.860000 418.320000 124.340000 ;
        RECT 417.120000 134.740000 418.320000 135.220000 ;
        RECT 462.120000 118.420000 463.320000 118.900000 ;
        RECT 462.120000 112.980000 463.320000 113.460000 ;
        RECT 462.120000 107.540000 463.320000 108.020000 ;
        RECT 462.120000 129.300000 463.320000 129.780000 ;
        RECT 462.120000 123.860000 463.320000 124.340000 ;
        RECT 462.120000 134.740000 463.320000 135.220000 ;
        RECT 507.120000 80.340000 508.320000 80.820000 ;
        RECT 507.120000 74.900000 508.320000 75.380000 ;
        RECT 507.120000 69.460000 508.320000 69.940000 ;
        RECT 507.120000 85.780000 508.320000 86.260000 ;
        RECT 507.120000 91.220000 508.320000 91.700000 ;
        RECT 507.120000 96.660000 508.320000 97.140000 ;
        RECT 507.120000 102.100000 508.320000 102.580000 ;
        RECT 543.400000 80.340000 544.600000 80.820000 ;
        RECT 543.400000 74.900000 544.600000 75.380000 ;
        RECT 543.400000 69.460000 544.600000 69.940000 ;
        RECT 543.400000 102.100000 544.600000 102.580000 ;
        RECT 543.400000 96.660000 544.600000 97.140000 ;
        RECT 543.400000 91.220000 544.600000 91.700000 ;
        RECT 543.400000 85.780000 544.600000 86.260000 ;
        RECT 507.120000 107.540000 508.320000 108.020000 ;
        RECT 507.120000 112.980000 508.320000 113.460000 ;
        RECT 507.120000 118.420000 508.320000 118.900000 ;
        RECT 507.120000 134.740000 508.320000 135.220000 ;
        RECT 507.120000 129.300000 508.320000 129.780000 ;
        RECT 507.120000 123.860000 508.320000 124.340000 ;
        RECT 543.400000 118.420000 544.600000 118.900000 ;
        RECT 543.400000 112.980000 544.600000 113.460000 ;
        RECT 543.400000 107.540000 544.600000 108.020000 ;
        RECT 543.400000 134.740000 544.600000 135.220000 ;
        RECT 543.400000 129.300000 544.600000 129.780000 ;
        RECT 543.400000 123.860000 544.600000 124.340000 ;
        RECT 282.120000 145.620000 283.320000 146.100000 ;
        RECT 282.120000 140.180000 283.320000 140.660000 ;
        RECT 282.120000 151.060000 283.320000 151.540000 ;
        RECT 282.120000 167.380000 283.320000 167.860000 ;
        RECT 282.120000 156.500000 283.320000 156.980000 ;
        RECT 282.120000 161.940000 283.320000 162.420000 ;
        RECT 327.120000 145.620000 328.320000 146.100000 ;
        RECT 327.120000 140.180000 328.320000 140.660000 ;
        RECT 327.120000 151.060000 328.320000 151.540000 ;
        RECT 327.120000 156.500000 328.320000 156.980000 ;
        RECT 327.120000 161.940000 328.320000 162.420000 ;
        RECT 327.120000 167.380000 328.320000 167.860000 ;
        RECT 282.120000 183.700000 283.320000 184.180000 ;
        RECT 282.120000 178.260000 283.320000 178.740000 ;
        RECT 282.120000 172.820000 283.320000 173.300000 ;
        RECT 282.120000 194.580000 283.320000 195.060000 ;
        RECT 282.120000 189.140000 283.320000 189.620000 ;
        RECT 282.120000 200.020000 283.320000 200.500000 ;
        RECT 282.120000 205.460000 283.320000 205.940000 ;
        RECT 327.120000 183.700000 328.320000 184.180000 ;
        RECT 327.120000 178.260000 328.320000 178.740000 ;
        RECT 327.120000 172.820000 328.320000 173.300000 ;
        RECT 327.120000 194.580000 328.320000 195.060000 ;
        RECT 327.120000 189.140000 328.320000 189.620000 ;
        RECT 327.120000 200.020000 328.320000 200.500000 ;
        RECT 327.120000 205.460000 328.320000 205.940000 ;
        RECT 372.120000 145.620000 373.320000 146.100000 ;
        RECT 372.120000 140.180000 373.320000 140.660000 ;
        RECT 372.120000 151.060000 373.320000 151.540000 ;
        RECT 372.120000 156.500000 373.320000 156.980000 ;
        RECT 372.120000 161.940000 373.320000 162.420000 ;
        RECT 372.120000 167.380000 373.320000 167.860000 ;
        RECT 372.120000 172.820000 373.320000 173.300000 ;
        RECT 372.120000 178.260000 373.320000 178.740000 ;
        RECT 372.120000 183.700000 373.320000 184.180000 ;
        RECT 372.120000 205.460000 373.320000 205.940000 ;
        RECT 372.120000 200.020000 373.320000 200.500000 ;
        RECT 372.120000 194.580000 373.320000 195.060000 ;
        RECT 372.120000 189.140000 373.320000 189.620000 ;
        RECT 282.120000 221.780000 283.320000 222.260000 ;
        RECT 282.120000 216.340000 283.320000 216.820000 ;
        RECT 282.120000 210.900000 283.320000 211.380000 ;
        RECT 282.120000 238.100000 283.320000 238.580000 ;
        RECT 282.120000 227.220000 283.320000 227.700000 ;
        RECT 282.120000 232.660000 283.320000 233.140000 ;
        RECT 327.120000 221.780000 328.320000 222.260000 ;
        RECT 327.120000 216.340000 328.320000 216.820000 ;
        RECT 327.120000 210.900000 328.320000 211.380000 ;
        RECT 327.120000 227.220000 328.320000 227.700000 ;
        RECT 327.120000 232.660000 328.320000 233.140000 ;
        RECT 327.120000 238.100000 328.320000 238.580000 ;
        RECT 282.120000 254.420000 283.320000 254.900000 ;
        RECT 282.120000 248.980000 283.320000 249.460000 ;
        RECT 282.120000 243.540000 283.320000 244.020000 ;
        RECT 282.120000 265.300000 283.320000 265.780000 ;
        RECT 282.120000 259.860000 283.320000 260.340000 ;
        RECT 282.120000 270.740000 283.320000 271.220000 ;
        RECT 327.120000 254.420000 328.320000 254.900000 ;
        RECT 327.120000 248.980000 328.320000 249.460000 ;
        RECT 327.120000 243.540000 328.320000 244.020000 ;
        RECT 327.120000 265.300000 328.320000 265.780000 ;
        RECT 327.120000 259.860000 328.320000 260.340000 ;
        RECT 327.120000 270.740000 328.320000 271.220000 ;
        RECT 372.120000 221.780000 373.320000 222.260000 ;
        RECT 372.120000 216.340000 373.320000 216.820000 ;
        RECT 372.120000 210.900000 373.320000 211.380000 ;
        RECT 372.120000 227.220000 373.320000 227.700000 ;
        RECT 372.120000 232.660000 373.320000 233.140000 ;
        RECT 372.120000 238.100000 373.320000 238.580000 ;
        RECT 372.120000 243.540000 373.320000 244.020000 ;
        RECT 372.120000 248.980000 373.320000 249.460000 ;
        RECT 372.120000 254.420000 373.320000 254.900000 ;
        RECT 372.120000 270.740000 373.320000 271.220000 ;
        RECT 372.120000 265.300000 373.320000 265.780000 ;
        RECT 372.120000 259.860000 373.320000 260.340000 ;
        RECT 417.120000 145.620000 418.320000 146.100000 ;
        RECT 417.120000 140.180000 418.320000 140.660000 ;
        RECT 417.120000 151.060000 418.320000 151.540000 ;
        RECT 417.120000 167.380000 418.320000 167.860000 ;
        RECT 417.120000 156.500000 418.320000 156.980000 ;
        RECT 417.120000 161.940000 418.320000 162.420000 ;
        RECT 462.120000 140.180000 463.320000 140.660000 ;
        RECT 462.120000 145.620000 463.320000 146.100000 ;
        RECT 462.120000 151.060000 463.320000 151.540000 ;
        RECT 462.120000 156.500000 463.320000 156.980000 ;
        RECT 462.120000 161.940000 463.320000 162.420000 ;
        RECT 462.120000 167.380000 463.320000 167.860000 ;
        RECT 417.120000 183.700000 418.320000 184.180000 ;
        RECT 417.120000 178.260000 418.320000 178.740000 ;
        RECT 417.120000 172.820000 418.320000 173.300000 ;
        RECT 417.120000 194.580000 418.320000 195.060000 ;
        RECT 417.120000 189.140000 418.320000 189.620000 ;
        RECT 417.120000 200.020000 418.320000 200.500000 ;
        RECT 417.120000 205.460000 418.320000 205.940000 ;
        RECT 462.120000 183.700000 463.320000 184.180000 ;
        RECT 462.120000 178.260000 463.320000 178.740000 ;
        RECT 462.120000 172.820000 463.320000 173.300000 ;
        RECT 462.120000 194.580000 463.320000 195.060000 ;
        RECT 462.120000 189.140000 463.320000 189.620000 ;
        RECT 462.120000 200.020000 463.320000 200.500000 ;
        RECT 462.120000 205.460000 463.320000 205.940000 ;
        RECT 507.120000 140.180000 508.320000 140.660000 ;
        RECT 507.120000 145.620000 508.320000 146.100000 ;
        RECT 507.120000 151.060000 508.320000 151.540000 ;
        RECT 507.120000 156.500000 508.320000 156.980000 ;
        RECT 507.120000 161.940000 508.320000 162.420000 ;
        RECT 507.120000 167.380000 508.320000 167.860000 ;
        RECT 543.400000 151.060000 544.600000 151.540000 ;
        RECT 543.400000 145.620000 544.600000 146.100000 ;
        RECT 543.400000 140.180000 544.600000 140.660000 ;
        RECT 543.400000 167.380000 544.600000 167.860000 ;
        RECT 543.400000 161.940000 544.600000 162.420000 ;
        RECT 543.400000 156.500000 544.600000 156.980000 ;
        RECT 507.120000 172.820000 508.320000 173.300000 ;
        RECT 507.120000 178.260000 508.320000 178.740000 ;
        RECT 507.120000 183.700000 508.320000 184.180000 ;
        RECT 507.120000 205.460000 508.320000 205.940000 ;
        RECT 507.120000 200.020000 508.320000 200.500000 ;
        RECT 507.120000 194.580000 508.320000 195.060000 ;
        RECT 507.120000 189.140000 508.320000 189.620000 ;
        RECT 543.400000 183.700000 544.600000 184.180000 ;
        RECT 543.400000 178.260000 544.600000 178.740000 ;
        RECT 543.400000 172.820000 544.600000 173.300000 ;
        RECT 543.400000 205.460000 544.600000 205.940000 ;
        RECT 543.400000 200.020000 544.600000 200.500000 ;
        RECT 543.400000 194.580000 544.600000 195.060000 ;
        RECT 543.400000 189.140000 544.600000 189.620000 ;
        RECT 417.120000 221.780000 418.320000 222.260000 ;
        RECT 417.120000 216.340000 418.320000 216.820000 ;
        RECT 417.120000 210.900000 418.320000 211.380000 ;
        RECT 417.120000 238.100000 418.320000 238.580000 ;
        RECT 417.120000 227.220000 418.320000 227.700000 ;
        RECT 417.120000 232.660000 418.320000 233.140000 ;
        RECT 462.120000 221.780000 463.320000 222.260000 ;
        RECT 462.120000 216.340000 463.320000 216.820000 ;
        RECT 462.120000 210.900000 463.320000 211.380000 ;
        RECT 462.120000 227.220000 463.320000 227.700000 ;
        RECT 462.120000 232.660000 463.320000 233.140000 ;
        RECT 462.120000 238.100000 463.320000 238.580000 ;
        RECT 417.120000 254.420000 418.320000 254.900000 ;
        RECT 417.120000 248.980000 418.320000 249.460000 ;
        RECT 417.120000 243.540000 418.320000 244.020000 ;
        RECT 417.120000 265.300000 418.320000 265.780000 ;
        RECT 417.120000 259.860000 418.320000 260.340000 ;
        RECT 417.120000 270.740000 418.320000 271.220000 ;
        RECT 462.120000 254.420000 463.320000 254.900000 ;
        RECT 462.120000 248.980000 463.320000 249.460000 ;
        RECT 462.120000 243.540000 463.320000 244.020000 ;
        RECT 462.120000 265.300000 463.320000 265.780000 ;
        RECT 462.120000 259.860000 463.320000 260.340000 ;
        RECT 462.120000 270.740000 463.320000 271.220000 ;
        RECT 507.120000 221.780000 508.320000 222.260000 ;
        RECT 507.120000 216.340000 508.320000 216.820000 ;
        RECT 507.120000 210.900000 508.320000 211.380000 ;
        RECT 507.120000 227.220000 508.320000 227.700000 ;
        RECT 507.120000 232.660000 508.320000 233.140000 ;
        RECT 507.120000 238.100000 508.320000 238.580000 ;
        RECT 543.400000 221.780000 544.600000 222.260000 ;
        RECT 543.400000 216.340000 544.600000 216.820000 ;
        RECT 543.400000 210.900000 544.600000 211.380000 ;
        RECT 543.400000 238.100000 544.600000 238.580000 ;
        RECT 543.400000 232.660000 544.600000 233.140000 ;
        RECT 543.400000 227.220000 544.600000 227.700000 ;
        RECT 507.120000 243.540000 508.320000 244.020000 ;
        RECT 507.120000 248.980000 508.320000 249.460000 ;
        RECT 507.120000 254.420000 508.320000 254.900000 ;
        RECT 507.120000 270.740000 508.320000 271.220000 ;
        RECT 507.120000 265.300000 508.320000 265.780000 ;
        RECT 507.120000 259.860000 508.320000 260.340000 ;
        RECT 543.400000 254.420000 544.600000 254.900000 ;
        RECT 543.400000 248.980000 544.600000 249.460000 ;
        RECT 543.400000 243.540000 544.600000 244.020000 ;
        RECT 543.400000 270.740000 544.600000 271.220000 ;
        RECT 543.400000 265.300000 544.600000 265.780000 ;
        RECT 543.400000 259.860000 544.600000 260.340000 ;
        RECT 5.560000 412.180000 6.760000 412.660000 ;
        RECT 192.120000 412.180000 193.320000 412.660000 ;
        RECT 147.120000 412.180000 148.320000 412.660000 ;
        RECT 102.120000 412.180000 103.320000 412.660000 ;
        RECT 57.120000 412.180000 58.320000 412.660000 ;
        RECT 12.120000 412.180000 13.320000 412.660000 ;
        RECT 237.120000 412.180000 238.320000 412.660000 ;
        RECT 5.560000 308.820000 6.760000 309.300000 ;
        RECT 57.120000 308.820000 58.320000 309.300000 ;
        RECT 12.120000 308.820000 13.320000 309.300000 ;
        RECT 5.560000 276.180000 6.760000 276.660000 ;
        RECT 5.560000 281.620000 6.760000 282.100000 ;
        RECT 12.120000 281.620000 13.320000 282.100000 ;
        RECT 12.120000 276.180000 13.320000 276.660000 ;
        RECT 5.560000 287.060000 6.760000 287.540000 ;
        RECT 12.120000 287.060000 13.320000 287.540000 ;
        RECT 5.560000 292.500000 6.760000 292.980000 ;
        RECT 5.560000 297.940000 6.760000 298.420000 ;
        RECT 12.120000 292.500000 13.320000 292.980000 ;
        RECT 12.120000 297.940000 13.320000 298.420000 ;
        RECT 5.560000 303.380000 6.760000 303.860000 ;
        RECT 12.120000 303.380000 13.320000 303.860000 ;
        RECT 57.120000 281.620000 58.320000 282.100000 ;
        RECT 57.120000 276.180000 58.320000 276.660000 ;
        RECT 57.120000 287.060000 58.320000 287.540000 ;
        RECT 57.120000 292.500000 58.320000 292.980000 ;
        RECT 57.120000 297.940000 58.320000 298.420000 ;
        RECT 57.120000 303.380000 58.320000 303.860000 ;
        RECT 5.560000 314.260000 6.760000 314.740000 ;
        RECT 12.120000 314.260000 13.320000 314.740000 ;
        RECT 5.560000 319.700000 6.760000 320.180000 ;
        RECT 5.560000 325.140000 6.760000 325.620000 ;
        RECT 12.120000 325.140000 13.320000 325.620000 ;
        RECT 12.120000 319.700000 13.320000 320.180000 ;
        RECT 5.560000 330.580000 6.760000 331.060000 ;
        RECT 12.120000 330.580000 13.320000 331.060000 ;
        RECT 5.560000 336.020000 6.760000 336.500000 ;
        RECT 5.560000 341.460000 6.760000 341.940000 ;
        RECT 12.120000 336.020000 13.320000 336.500000 ;
        RECT 12.120000 341.460000 13.320000 341.940000 ;
        RECT 57.120000 325.140000 58.320000 325.620000 ;
        RECT 57.120000 319.700000 58.320000 320.180000 ;
        RECT 57.120000 314.260000 58.320000 314.740000 ;
        RECT 57.120000 336.020000 58.320000 336.500000 ;
        RECT 57.120000 330.580000 58.320000 331.060000 ;
        RECT 57.120000 341.460000 58.320000 341.940000 ;
        RECT 102.120000 308.820000 103.320000 309.300000 ;
        RECT 102.120000 281.620000 103.320000 282.100000 ;
        RECT 102.120000 276.180000 103.320000 276.660000 ;
        RECT 102.120000 287.060000 103.320000 287.540000 ;
        RECT 102.120000 292.500000 103.320000 292.980000 ;
        RECT 102.120000 297.940000 103.320000 298.420000 ;
        RECT 102.120000 303.380000 103.320000 303.860000 ;
        RECT 102.120000 341.460000 103.320000 341.940000 ;
        RECT 102.120000 336.020000 103.320000 336.500000 ;
        RECT 102.120000 330.580000 103.320000 331.060000 ;
        RECT 102.120000 314.260000 103.320000 314.740000 ;
        RECT 102.120000 319.700000 103.320000 320.180000 ;
        RECT 102.120000 325.140000 103.320000 325.620000 ;
        RECT 5.560000 346.900000 6.760000 347.380000 ;
        RECT 12.120000 346.900000 13.320000 347.380000 ;
        RECT 5.560000 352.340000 6.760000 352.820000 ;
        RECT 5.560000 357.780000 6.760000 358.260000 ;
        RECT 12.120000 357.780000 13.320000 358.260000 ;
        RECT 12.120000 352.340000 13.320000 352.820000 ;
        RECT 5.560000 363.220000 6.760000 363.700000 ;
        RECT 5.560000 368.660000 6.760000 369.140000 ;
        RECT 12.120000 363.220000 13.320000 363.700000 ;
        RECT 12.120000 368.660000 13.320000 369.140000 ;
        RECT 5.560000 374.100000 6.760000 374.580000 ;
        RECT 12.120000 374.100000 13.320000 374.580000 ;
        RECT 57.120000 357.780000 58.320000 358.260000 ;
        RECT 57.120000 352.340000 58.320000 352.820000 ;
        RECT 57.120000 346.900000 58.320000 347.380000 ;
        RECT 57.120000 363.220000 58.320000 363.700000 ;
        RECT 57.120000 368.660000 58.320000 369.140000 ;
        RECT 57.120000 374.100000 58.320000 374.580000 ;
        RECT 5.560000 379.540000 6.760000 380.020000 ;
        RECT 5.560000 384.980000 6.760000 385.460000 ;
        RECT 12.120000 384.980000 13.320000 385.460000 ;
        RECT 12.120000 379.540000 13.320000 380.020000 ;
        RECT 5.560000 390.420000 6.760000 390.900000 ;
        RECT 12.120000 390.420000 13.320000 390.900000 ;
        RECT 5.560000 395.860000 6.760000 396.340000 ;
        RECT 5.560000 401.300000 6.760000 401.780000 ;
        RECT 12.120000 401.300000 13.320000 401.780000 ;
        RECT 12.120000 395.860000 13.320000 396.340000 ;
        RECT 5.560000 406.740000 6.760000 407.220000 ;
        RECT 12.120000 406.740000 13.320000 407.220000 ;
        RECT 57.120000 390.420000 58.320000 390.900000 ;
        RECT 57.120000 384.980000 58.320000 385.460000 ;
        RECT 57.120000 379.540000 58.320000 380.020000 ;
        RECT 57.120000 401.300000 58.320000 401.780000 ;
        RECT 57.120000 395.860000 58.320000 396.340000 ;
        RECT 57.120000 406.740000 58.320000 407.220000 ;
        RECT 102.120000 357.780000 103.320000 358.260000 ;
        RECT 102.120000 352.340000 103.320000 352.820000 ;
        RECT 102.120000 346.900000 103.320000 347.380000 ;
        RECT 102.120000 363.220000 103.320000 363.700000 ;
        RECT 102.120000 368.660000 103.320000 369.140000 ;
        RECT 102.120000 374.100000 103.320000 374.580000 ;
        RECT 102.120000 406.740000 103.320000 407.220000 ;
        RECT 102.120000 401.300000 103.320000 401.780000 ;
        RECT 102.120000 379.540000 103.320000 380.020000 ;
        RECT 102.120000 384.980000 103.320000 385.460000 ;
        RECT 102.120000 390.420000 103.320000 390.900000 ;
        RECT 102.120000 395.860000 103.320000 396.340000 ;
        RECT 192.120000 308.820000 193.320000 309.300000 ;
        RECT 147.120000 308.820000 148.320000 309.300000 ;
        RECT 147.120000 276.180000 148.320000 276.660000 ;
        RECT 147.120000 281.620000 148.320000 282.100000 ;
        RECT 147.120000 287.060000 148.320000 287.540000 ;
        RECT 147.120000 303.380000 148.320000 303.860000 ;
        RECT 147.120000 292.500000 148.320000 292.980000 ;
        RECT 147.120000 297.940000 148.320000 298.420000 ;
        RECT 192.120000 276.180000 193.320000 276.660000 ;
        RECT 192.120000 281.620000 193.320000 282.100000 ;
        RECT 192.120000 287.060000 193.320000 287.540000 ;
        RECT 192.120000 292.500000 193.320000 292.980000 ;
        RECT 192.120000 297.940000 193.320000 298.420000 ;
        RECT 192.120000 303.380000 193.320000 303.860000 ;
        RECT 147.120000 325.140000 148.320000 325.620000 ;
        RECT 147.120000 319.700000 148.320000 320.180000 ;
        RECT 147.120000 314.260000 148.320000 314.740000 ;
        RECT 147.120000 336.020000 148.320000 336.500000 ;
        RECT 147.120000 330.580000 148.320000 331.060000 ;
        RECT 147.120000 341.460000 148.320000 341.940000 ;
        RECT 192.120000 325.140000 193.320000 325.620000 ;
        RECT 192.120000 319.700000 193.320000 320.180000 ;
        RECT 192.120000 314.260000 193.320000 314.740000 ;
        RECT 192.120000 336.020000 193.320000 336.500000 ;
        RECT 192.120000 330.580000 193.320000 331.060000 ;
        RECT 192.120000 341.460000 193.320000 341.940000 ;
        RECT 237.120000 308.820000 238.320000 309.300000 ;
        RECT 237.120000 281.620000 238.320000 282.100000 ;
        RECT 237.120000 276.180000 238.320000 276.660000 ;
        RECT 237.120000 287.060000 238.320000 287.540000 ;
        RECT 237.120000 292.500000 238.320000 292.980000 ;
        RECT 237.120000 297.940000 238.320000 298.420000 ;
        RECT 237.120000 303.380000 238.320000 303.860000 ;
        RECT 237.120000 314.260000 238.320000 314.740000 ;
        RECT 237.120000 319.700000 238.320000 320.180000 ;
        RECT 237.120000 325.140000 238.320000 325.620000 ;
        RECT 237.120000 341.460000 238.320000 341.940000 ;
        RECT 237.120000 336.020000 238.320000 336.500000 ;
        RECT 237.120000 330.580000 238.320000 331.060000 ;
        RECT 147.120000 357.780000 148.320000 358.260000 ;
        RECT 147.120000 352.340000 148.320000 352.820000 ;
        RECT 147.120000 346.900000 148.320000 347.380000 ;
        RECT 147.120000 374.100000 148.320000 374.580000 ;
        RECT 147.120000 363.220000 148.320000 363.700000 ;
        RECT 147.120000 368.660000 148.320000 369.140000 ;
        RECT 192.120000 357.780000 193.320000 358.260000 ;
        RECT 192.120000 352.340000 193.320000 352.820000 ;
        RECT 192.120000 346.900000 193.320000 347.380000 ;
        RECT 192.120000 363.220000 193.320000 363.700000 ;
        RECT 192.120000 368.660000 193.320000 369.140000 ;
        RECT 192.120000 374.100000 193.320000 374.580000 ;
        RECT 147.120000 390.420000 148.320000 390.900000 ;
        RECT 147.120000 384.980000 148.320000 385.460000 ;
        RECT 147.120000 379.540000 148.320000 380.020000 ;
        RECT 147.120000 401.300000 148.320000 401.780000 ;
        RECT 147.120000 395.860000 148.320000 396.340000 ;
        RECT 147.120000 406.740000 148.320000 407.220000 ;
        RECT 192.120000 390.420000 193.320000 390.900000 ;
        RECT 192.120000 384.980000 193.320000 385.460000 ;
        RECT 192.120000 379.540000 193.320000 380.020000 ;
        RECT 192.120000 401.300000 193.320000 401.780000 ;
        RECT 192.120000 395.860000 193.320000 396.340000 ;
        RECT 192.120000 406.740000 193.320000 407.220000 ;
        RECT 237.120000 357.780000 238.320000 358.260000 ;
        RECT 237.120000 352.340000 238.320000 352.820000 ;
        RECT 237.120000 346.900000 238.320000 347.380000 ;
        RECT 237.120000 363.220000 238.320000 363.700000 ;
        RECT 237.120000 368.660000 238.320000 369.140000 ;
        RECT 237.120000 374.100000 238.320000 374.580000 ;
        RECT 237.120000 379.540000 238.320000 380.020000 ;
        RECT 237.120000 384.980000 238.320000 385.460000 ;
        RECT 237.120000 390.420000 238.320000 390.900000 ;
        RECT 237.120000 406.740000 238.320000 407.220000 ;
        RECT 237.120000 401.300000 238.320000 401.780000 ;
        RECT 237.120000 395.860000 238.320000 396.340000 ;
        RECT 5.560000 417.620000 6.760000 418.100000 ;
        RECT 12.120000 417.620000 13.320000 418.100000 ;
        RECT 5.560000 423.060000 6.760000 423.540000 ;
        RECT 5.560000 428.500000 6.760000 428.980000 ;
        RECT 12.120000 423.060000 13.320000 423.540000 ;
        RECT 12.120000 428.500000 13.320000 428.980000 ;
        RECT 5.560000 433.940000 6.760000 434.420000 ;
        RECT 12.120000 433.940000 13.320000 434.420000 ;
        RECT 5.560000 439.380000 6.760000 439.860000 ;
        RECT 5.560000 444.820000 6.760000 445.300000 ;
        RECT 12.120000 444.820000 13.320000 445.300000 ;
        RECT 12.120000 439.380000 13.320000 439.860000 ;
        RECT 57.120000 417.620000 58.320000 418.100000 ;
        RECT 57.120000 423.060000 58.320000 423.540000 ;
        RECT 57.120000 428.500000 58.320000 428.980000 ;
        RECT 57.120000 433.940000 58.320000 434.420000 ;
        RECT 57.120000 439.380000 58.320000 439.860000 ;
        RECT 57.120000 444.820000 58.320000 445.300000 ;
        RECT 5.560000 450.260000 6.760000 450.740000 ;
        RECT 12.120000 450.260000 13.320000 450.740000 ;
        RECT 5.560000 455.700000 6.760000 456.180000 ;
        RECT 5.560000 461.140000 6.760000 461.620000 ;
        RECT 12.120000 461.140000 13.320000 461.620000 ;
        RECT 12.120000 455.700000 13.320000 456.180000 ;
        RECT 5.560000 466.580000 6.760000 467.060000 ;
        RECT 5.560000 472.020000 6.760000 472.500000 ;
        RECT 12.120000 472.020000 13.320000 472.500000 ;
        RECT 12.120000 466.580000 13.320000 467.060000 ;
        RECT 5.560000 477.460000 6.760000 477.940000 ;
        RECT 12.120000 477.460000 13.320000 477.940000 ;
        RECT 57.120000 461.140000 58.320000 461.620000 ;
        RECT 57.120000 455.700000 58.320000 456.180000 ;
        RECT 57.120000 450.260000 58.320000 450.740000 ;
        RECT 57.120000 472.020000 58.320000 472.500000 ;
        RECT 57.120000 466.580000 58.320000 467.060000 ;
        RECT 57.120000 477.460000 58.320000 477.940000 ;
        RECT 102.120000 428.500000 103.320000 428.980000 ;
        RECT 102.120000 417.620000 103.320000 418.100000 ;
        RECT 102.120000 423.060000 103.320000 423.540000 ;
        RECT 102.120000 433.940000 103.320000 434.420000 ;
        RECT 102.120000 439.380000 103.320000 439.860000 ;
        RECT 102.120000 444.820000 103.320000 445.300000 ;
        RECT 102.120000 477.460000 103.320000 477.940000 ;
        RECT 102.120000 472.020000 103.320000 472.500000 ;
        RECT 102.120000 450.260000 103.320000 450.740000 ;
        RECT 102.120000 455.700000 103.320000 456.180000 ;
        RECT 102.120000 461.140000 103.320000 461.620000 ;
        RECT 102.120000 466.580000 103.320000 467.060000 ;
        RECT 5.560000 515.540000 6.760000 516.020000 ;
        RECT 57.120000 515.540000 58.320000 516.020000 ;
        RECT 12.120000 515.540000 13.320000 516.020000 ;
        RECT 5.560000 482.900000 6.760000 483.380000 ;
        RECT 5.560000 488.340000 6.760000 488.820000 ;
        RECT 12.120000 488.340000 13.320000 488.820000 ;
        RECT 12.120000 482.900000 13.320000 483.380000 ;
        RECT 5.560000 493.780000 6.760000 494.260000 ;
        RECT 12.120000 493.780000 13.320000 494.260000 ;
        RECT 5.560000 499.220000 6.760000 499.700000 ;
        RECT 5.560000 504.660000 6.760000 505.140000 ;
        RECT 12.120000 504.660000 13.320000 505.140000 ;
        RECT 12.120000 499.220000 13.320000 499.700000 ;
        RECT 5.560000 510.100000 6.760000 510.580000 ;
        RECT 12.120000 510.100000 13.320000 510.580000 ;
        RECT 57.120000 493.780000 58.320000 494.260000 ;
        RECT 57.120000 488.340000 58.320000 488.820000 ;
        RECT 57.120000 482.900000 58.320000 483.380000 ;
        RECT 57.120000 504.660000 58.320000 505.140000 ;
        RECT 57.120000 499.220000 58.320000 499.700000 ;
        RECT 57.120000 510.100000 58.320000 510.580000 ;
        RECT 5.560000 520.980000 6.760000 521.460000 ;
        RECT 12.120000 520.980000 13.320000 521.460000 ;
        RECT 5.560000 526.420000 6.760000 526.900000 ;
        RECT 5.560000 531.860000 6.760000 532.340000 ;
        RECT 12.120000 531.860000 13.320000 532.340000 ;
        RECT 12.120000 526.420000 13.320000 526.900000 ;
        RECT 12.120000 537.300000 13.320000 537.780000 ;
        RECT 5.560000 537.300000 6.760000 537.780000 ;
        RECT 57.120000 520.980000 58.320000 521.460000 ;
        RECT 57.120000 526.420000 58.320000 526.900000 ;
        RECT 57.120000 531.860000 58.320000 532.340000 ;
        RECT 57.120000 537.300000 58.320000 537.780000 ;
        RECT 102.120000 515.540000 103.320000 516.020000 ;
        RECT 102.120000 488.340000 103.320000 488.820000 ;
        RECT 102.120000 482.900000 103.320000 483.380000 ;
        RECT 102.120000 493.780000 103.320000 494.260000 ;
        RECT 102.120000 499.220000 103.320000 499.700000 ;
        RECT 102.120000 504.660000 103.320000 505.140000 ;
        RECT 102.120000 510.100000 103.320000 510.580000 ;
        RECT 102.120000 537.300000 103.320000 537.780000 ;
        RECT 102.120000 520.980000 103.320000 521.460000 ;
        RECT 102.120000 526.420000 103.320000 526.900000 ;
        RECT 102.120000 531.860000 103.320000 532.340000 ;
        RECT 147.120000 417.620000 148.320000 418.100000 ;
        RECT 147.120000 423.060000 148.320000 423.540000 ;
        RECT 147.120000 428.500000 148.320000 428.980000 ;
        RECT 147.120000 444.820000 148.320000 445.300000 ;
        RECT 147.120000 433.940000 148.320000 434.420000 ;
        RECT 147.120000 439.380000 148.320000 439.860000 ;
        RECT 192.120000 428.500000 193.320000 428.980000 ;
        RECT 192.120000 417.620000 193.320000 418.100000 ;
        RECT 192.120000 423.060000 193.320000 423.540000 ;
        RECT 192.120000 433.940000 193.320000 434.420000 ;
        RECT 192.120000 439.380000 193.320000 439.860000 ;
        RECT 192.120000 444.820000 193.320000 445.300000 ;
        RECT 147.120000 461.140000 148.320000 461.620000 ;
        RECT 147.120000 455.700000 148.320000 456.180000 ;
        RECT 147.120000 450.260000 148.320000 450.740000 ;
        RECT 147.120000 472.020000 148.320000 472.500000 ;
        RECT 147.120000 466.580000 148.320000 467.060000 ;
        RECT 147.120000 477.460000 148.320000 477.940000 ;
        RECT 192.120000 461.140000 193.320000 461.620000 ;
        RECT 192.120000 455.700000 193.320000 456.180000 ;
        RECT 192.120000 450.260000 193.320000 450.740000 ;
        RECT 192.120000 472.020000 193.320000 472.500000 ;
        RECT 192.120000 466.580000 193.320000 467.060000 ;
        RECT 192.120000 477.460000 193.320000 477.940000 ;
        RECT 237.120000 417.620000 238.320000 418.100000 ;
        RECT 237.120000 423.060000 238.320000 423.540000 ;
        RECT 237.120000 428.500000 238.320000 428.980000 ;
        RECT 237.120000 433.940000 238.320000 434.420000 ;
        RECT 237.120000 439.380000 238.320000 439.860000 ;
        RECT 237.120000 444.820000 238.320000 445.300000 ;
        RECT 237.120000 450.260000 238.320000 450.740000 ;
        RECT 237.120000 455.700000 238.320000 456.180000 ;
        RECT 237.120000 461.140000 238.320000 461.620000 ;
        RECT 237.120000 477.460000 238.320000 477.940000 ;
        RECT 237.120000 472.020000 238.320000 472.500000 ;
        RECT 237.120000 466.580000 238.320000 467.060000 ;
        RECT 192.120000 515.540000 193.320000 516.020000 ;
        RECT 147.120000 515.540000 148.320000 516.020000 ;
        RECT 147.120000 493.780000 148.320000 494.260000 ;
        RECT 147.120000 488.340000 148.320000 488.820000 ;
        RECT 147.120000 482.900000 148.320000 483.380000 ;
        RECT 147.120000 499.220000 148.320000 499.700000 ;
        RECT 147.120000 504.660000 148.320000 505.140000 ;
        RECT 147.120000 510.100000 148.320000 510.580000 ;
        RECT 192.120000 488.340000 193.320000 488.820000 ;
        RECT 192.120000 482.900000 193.320000 483.380000 ;
        RECT 192.120000 493.780000 193.320000 494.260000 ;
        RECT 192.120000 504.660000 193.320000 505.140000 ;
        RECT 192.120000 499.220000 193.320000 499.700000 ;
        RECT 192.120000 510.100000 193.320000 510.580000 ;
        RECT 147.120000 520.980000 148.320000 521.460000 ;
        RECT 147.120000 526.420000 148.320000 526.900000 ;
        RECT 147.120000 531.860000 148.320000 532.340000 ;
        RECT 147.120000 537.300000 148.320000 537.780000 ;
        RECT 192.120000 520.980000 193.320000 521.460000 ;
        RECT 192.120000 526.420000 193.320000 526.900000 ;
        RECT 192.120000 531.860000 193.320000 532.340000 ;
        RECT 192.120000 537.300000 193.320000 537.780000 ;
        RECT 237.120000 515.540000 238.320000 516.020000 ;
        RECT 237.120000 493.780000 238.320000 494.260000 ;
        RECT 237.120000 488.340000 238.320000 488.820000 ;
        RECT 237.120000 482.900000 238.320000 483.380000 ;
        RECT 237.120000 499.220000 238.320000 499.700000 ;
        RECT 237.120000 504.660000 238.320000 505.140000 ;
        RECT 237.120000 510.100000 238.320000 510.580000 ;
        RECT 237.120000 537.300000 238.320000 537.780000 ;
        RECT 237.120000 520.980000 238.320000 521.460000 ;
        RECT 237.120000 526.420000 238.320000 526.900000 ;
        RECT 237.120000 531.860000 238.320000 532.340000 ;
        RECT 543.400000 412.180000 544.600000 412.660000 ;
        RECT 507.120000 412.180000 508.320000 412.660000 ;
        RECT 462.120000 412.180000 463.320000 412.660000 ;
        RECT 417.120000 412.180000 418.320000 412.660000 ;
        RECT 372.120000 412.180000 373.320000 412.660000 ;
        RECT 327.120000 412.180000 328.320000 412.660000 ;
        RECT 282.120000 412.180000 283.320000 412.660000 ;
        RECT 327.120000 308.820000 328.320000 309.300000 ;
        RECT 282.120000 308.820000 283.320000 309.300000 ;
        RECT 282.120000 281.620000 283.320000 282.100000 ;
        RECT 282.120000 276.180000 283.320000 276.660000 ;
        RECT 282.120000 287.060000 283.320000 287.540000 ;
        RECT 282.120000 303.380000 283.320000 303.860000 ;
        RECT 282.120000 292.500000 283.320000 292.980000 ;
        RECT 282.120000 297.940000 283.320000 298.420000 ;
        RECT 327.120000 281.620000 328.320000 282.100000 ;
        RECT 327.120000 276.180000 328.320000 276.660000 ;
        RECT 327.120000 287.060000 328.320000 287.540000 ;
        RECT 327.120000 292.500000 328.320000 292.980000 ;
        RECT 327.120000 297.940000 328.320000 298.420000 ;
        RECT 327.120000 303.380000 328.320000 303.860000 ;
        RECT 282.120000 325.140000 283.320000 325.620000 ;
        RECT 282.120000 319.700000 283.320000 320.180000 ;
        RECT 282.120000 314.260000 283.320000 314.740000 ;
        RECT 282.120000 336.020000 283.320000 336.500000 ;
        RECT 282.120000 330.580000 283.320000 331.060000 ;
        RECT 282.120000 341.460000 283.320000 341.940000 ;
        RECT 327.120000 325.140000 328.320000 325.620000 ;
        RECT 327.120000 319.700000 328.320000 320.180000 ;
        RECT 327.120000 314.260000 328.320000 314.740000 ;
        RECT 327.120000 336.020000 328.320000 336.500000 ;
        RECT 327.120000 330.580000 328.320000 331.060000 ;
        RECT 327.120000 341.460000 328.320000 341.940000 ;
        RECT 372.120000 308.820000 373.320000 309.300000 ;
        RECT 372.120000 281.620000 373.320000 282.100000 ;
        RECT 372.120000 276.180000 373.320000 276.660000 ;
        RECT 372.120000 287.060000 373.320000 287.540000 ;
        RECT 372.120000 292.500000 373.320000 292.980000 ;
        RECT 372.120000 297.940000 373.320000 298.420000 ;
        RECT 372.120000 303.380000 373.320000 303.860000 ;
        RECT 372.120000 314.260000 373.320000 314.740000 ;
        RECT 372.120000 319.700000 373.320000 320.180000 ;
        RECT 372.120000 325.140000 373.320000 325.620000 ;
        RECT 372.120000 341.460000 373.320000 341.940000 ;
        RECT 372.120000 336.020000 373.320000 336.500000 ;
        RECT 372.120000 330.580000 373.320000 331.060000 ;
        RECT 282.120000 357.780000 283.320000 358.260000 ;
        RECT 282.120000 352.340000 283.320000 352.820000 ;
        RECT 282.120000 346.900000 283.320000 347.380000 ;
        RECT 282.120000 374.100000 283.320000 374.580000 ;
        RECT 282.120000 363.220000 283.320000 363.700000 ;
        RECT 282.120000 368.660000 283.320000 369.140000 ;
        RECT 327.120000 357.780000 328.320000 358.260000 ;
        RECT 327.120000 352.340000 328.320000 352.820000 ;
        RECT 327.120000 346.900000 328.320000 347.380000 ;
        RECT 327.120000 363.220000 328.320000 363.700000 ;
        RECT 327.120000 368.660000 328.320000 369.140000 ;
        RECT 327.120000 374.100000 328.320000 374.580000 ;
        RECT 282.120000 390.420000 283.320000 390.900000 ;
        RECT 282.120000 384.980000 283.320000 385.460000 ;
        RECT 282.120000 379.540000 283.320000 380.020000 ;
        RECT 282.120000 401.300000 283.320000 401.780000 ;
        RECT 282.120000 395.860000 283.320000 396.340000 ;
        RECT 282.120000 406.740000 283.320000 407.220000 ;
        RECT 327.120000 390.420000 328.320000 390.900000 ;
        RECT 327.120000 384.980000 328.320000 385.460000 ;
        RECT 327.120000 379.540000 328.320000 380.020000 ;
        RECT 327.120000 401.300000 328.320000 401.780000 ;
        RECT 327.120000 395.860000 328.320000 396.340000 ;
        RECT 327.120000 406.740000 328.320000 407.220000 ;
        RECT 372.120000 357.780000 373.320000 358.260000 ;
        RECT 372.120000 352.340000 373.320000 352.820000 ;
        RECT 372.120000 346.900000 373.320000 347.380000 ;
        RECT 372.120000 363.220000 373.320000 363.700000 ;
        RECT 372.120000 368.660000 373.320000 369.140000 ;
        RECT 372.120000 374.100000 373.320000 374.580000 ;
        RECT 372.120000 379.540000 373.320000 380.020000 ;
        RECT 372.120000 384.980000 373.320000 385.460000 ;
        RECT 372.120000 390.420000 373.320000 390.900000 ;
        RECT 372.120000 406.740000 373.320000 407.220000 ;
        RECT 372.120000 401.300000 373.320000 401.780000 ;
        RECT 372.120000 395.860000 373.320000 396.340000 ;
        RECT 462.120000 308.820000 463.320000 309.300000 ;
        RECT 417.120000 308.820000 418.320000 309.300000 ;
        RECT 417.120000 281.620000 418.320000 282.100000 ;
        RECT 417.120000 276.180000 418.320000 276.660000 ;
        RECT 417.120000 287.060000 418.320000 287.540000 ;
        RECT 417.120000 303.380000 418.320000 303.860000 ;
        RECT 417.120000 292.500000 418.320000 292.980000 ;
        RECT 417.120000 297.940000 418.320000 298.420000 ;
        RECT 462.120000 276.180000 463.320000 276.660000 ;
        RECT 462.120000 281.620000 463.320000 282.100000 ;
        RECT 462.120000 287.060000 463.320000 287.540000 ;
        RECT 462.120000 292.500000 463.320000 292.980000 ;
        RECT 462.120000 297.940000 463.320000 298.420000 ;
        RECT 462.120000 303.380000 463.320000 303.860000 ;
        RECT 417.120000 325.140000 418.320000 325.620000 ;
        RECT 417.120000 319.700000 418.320000 320.180000 ;
        RECT 417.120000 314.260000 418.320000 314.740000 ;
        RECT 417.120000 336.020000 418.320000 336.500000 ;
        RECT 417.120000 330.580000 418.320000 331.060000 ;
        RECT 417.120000 341.460000 418.320000 341.940000 ;
        RECT 462.120000 325.140000 463.320000 325.620000 ;
        RECT 462.120000 319.700000 463.320000 320.180000 ;
        RECT 462.120000 314.260000 463.320000 314.740000 ;
        RECT 462.120000 336.020000 463.320000 336.500000 ;
        RECT 462.120000 330.580000 463.320000 331.060000 ;
        RECT 462.120000 341.460000 463.320000 341.940000 ;
        RECT 543.400000 308.820000 544.600000 309.300000 ;
        RECT 507.120000 308.820000 508.320000 309.300000 ;
        RECT 507.120000 276.180000 508.320000 276.660000 ;
        RECT 507.120000 281.620000 508.320000 282.100000 ;
        RECT 507.120000 287.060000 508.320000 287.540000 ;
        RECT 507.120000 292.500000 508.320000 292.980000 ;
        RECT 507.120000 297.940000 508.320000 298.420000 ;
        RECT 507.120000 303.380000 508.320000 303.860000 ;
        RECT 543.400000 287.060000 544.600000 287.540000 ;
        RECT 543.400000 281.620000 544.600000 282.100000 ;
        RECT 543.400000 276.180000 544.600000 276.660000 ;
        RECT 543.400000 303.380000 544.600000 303.860000 ;
        RECT 543.400000 297.940000 544.600000 298.420000 ;
        RECT 543.400000 292.500000 544.600000 292.980000 ;
        RECT 507.120000 314.260000 508.320000 314.740000 ;
        RECT 507.120000 319.700000 508.320000 320.180000 ;
        RECT 507.120000 325.140000 508.320000 325.620000 ;
        RECT 507.120000 341.460000 508.320000 341.940000 ;
        RECT 507.120000 336.020000 508.320000 336.500000 ;
        RECT 507.120000 330.580000 508.320000 331.060000 ;
        RECT 543.400000 325.140000 544.600000 325.620000 ;
        RECT 543.400000 319.700000 544.600000 320.180000 ;
        RECT 543.400000 314.260000 544.600000 314.740000 ;
        RECT 543.400000 341.460000 544.600000 341.940000 ;
        RECT 543.400000 336.020000 544.600000 336.500000 ;
        RECT 543.400000 330.580000 544.600000 331.060000 ;
        RECT 417.120000 357.780000 418.320000 358.260000 ;
        RECT 417.120000 352.340000 418.320000 352.820000 ;
        RECT 417.120000 346.900000 418.320000 347.380000 ;
        RECT 417.120000 374.100000 418.320000 374.580000 ;
        RECT 417.120000 363.220000 418.320000 363.700000 ;
        RECT 417.120000 368.660000 418.320000 369.140000 ;
        RECT 462.120000 357.780000 463.320000 358.260000 ;
        RECT 462.120000 352.340000 463.320000 352.820000 ;
        RECT 462.120000 346.900000 463.320000 347.380000 ;
        RECT 462.120000 363.220000 463.320000 363.700000 ;
        RECT 462.120000 368.660000 463.320000 369.140000 ;
        RECT 462.120000 374.100000 463.320000 374.580000 ;
        RECT 417.120000 390.420000 418.320000 390.900000 ;
        RECT 417.120000 384.980000 418.320000 385.460000 ;
        RECT 417.120000 379.540000 418.320000 380.020000 ;
        RECT 417.120000 401.300000 418.320000 401.780000 ;
        RECT 417.120000 395.860000 418.320000 396.340000 ;
        RECT 417.120000 406.740000 418.320000 407.220000 ;
        RECT 462.120000 390.420000 463.320000 390.900000 ;
        RECT 462.120000 384.980000 463.320000 385.460000 ;
        RECT 462.120000 379.540000 463.320000 380.020000 ;
        RECT 462.120000 401.300000 463.320000 401.780000 ;
        RECT 462.120000 395.860000 463.320000 396.340000 ;
        RECT 462.120000 406.740000 463.320000 407.220000 ;
        RECT 507.120000 357.780000 508.320000 358.260000 ;
        RECT 507.120000 352.340000 508.320000 352.820000 ;
        RECT 507.120000 346.900000 508.320000 347.380000 ;
        RECT 507.120000 363.220000 508.320000 363.700000 ;
        RECT 507.120000 368.660000 508.320000 369.140000 ;
        RECT 507.120000 374.100000 508.320000 374.580000 ;
        RECT 543.400000 357.780000 544.600000 358.260000 ;
        RECT 543.400000 352.340000 544.600000 352.820000 ;
        RECT 543.400000 346.900000 544.600000 347.380000 ;
        RECT 543.400000 374.100000 544.600000 374.580000 ;
        RECT 543.400000 368.660000 544.600000 369.140000 ;
        RECT 543.400000 363.220000 544.600000 363.700000 ;
        RECT 507.120000 379.540000 508.320000 380.020000 ;
        RECT 507.120000 384.980000 508.320000 385.460000 ;
        RECT 507.120000 390.420000 508.320000 390.900000 ;
        RECT 507.120000 406.740000 508.320000 407.220000 ;
        RECT 507.120000 401.300000 508.320000 401.780000 ;
        RECT 507.120000 395.860000 508.320000 396.340000 ;
        RECT 543.400000 390.420000 544.600000 390.900000 ;
        RECT 543.400000 384.980000 544.600000 385.460000 ;
        RECT 543.400000 379.540000 544.600000 380.020000 ;
        RECT 543.400000 406.740000 544.600000 407.220000 ;
        RECT 543.400000 401.300000 544.600000 401.780000 ;
        RECT 543.400000 395.860000 544.600000 396.340000 ;
        RECT 282.120000 417.620000 283.320000 418.100000 ;
        RECT 282.120000 423.060000 283.320000 423.540000 ;
        RECT 282.120000 428.500000 283.320000 428.980000 ;
        RECT 282.120000 444.820000 283.320000 445.300000 ;
        RECT 282.120000 433.940000 283.320000 434.420000 ;
        RECT 282.120000 439.380000 283.320000 439.860000 ;
        RECT 327.120000 417.620000 328.320000 418.100000 ;
        RECT 327.120000 423.060000 328.320000 423.540000 ;
        RECT 327.120000 428.500000 328.320000 428.980000 ;
        RECT 327.120000 433.940000 328.320000 434.420000 ;
        RECT 327.120000 439.380000 328.320000 439.860000 ;
        RECT 327.120000 444.820000 328.320000 445.300000 ;
        RECT 282.120000 461.140000 283.320000 461.620000 ;
        RECT 282.120000 455.700000 283.320000 456.180000 ;
        RECT 282.120000 450.260000 283.320000 450.740000 ;
        RECT 282.120000 472.020000 283.320000 472.500000 ;
        RECT 282.120000 466.580000 283.320000 467.060000 ;
        RECT 282.120000 477.460000 283.320000 477.940000 ;
        RECT 327.120000 461.140000 328.320000 461.620000 ;
        RECT 327.120000 455.700000 328.320000 456.180000 ;
        RECT 327.120000 450.260000 328.320000 450.740000 ;
        RECT 327.120000 472.020000 328.320000 472.500000 ;
        RECT 327.120000 466.580000 328.320000 467.060000 ;
        RECT 327.120000 477.460000 328.320000 477.940000 ;
        RECT 372.120000 428.500000 373.320000 428.980000 ;
        RECT 372.120000 417.620000 373.320000 418.100000 ;
        RECT 372.120000 423.060000 373.320000 423.540000 ;
        RECT 372.120000 433.940000 373.320000 434.420000 ;
        RECT 372.120000 439.380000 373.320000 439.860000 ;
        RECT 372.120000 444.820000 373.320000 445.300000 ;
        RECT 372.120000 450.260000 373.320000 450.740000 ;
        RECT 372.120000 455.700000 373.320000 456.180000 ;
        RECT 372.120000 461.140000 373.320000 461.620000 ;
        RECT 372.120000 477.460000 373.320000 477.940000 ;
        RECT 372.120000 472.020000 373.320000 472.500000 ;
        RECT 372.120000 466.580000 373.320000 467.060000 ;
        RECT 327.120000 515.540000 328.320000 516.020000 ;
        RECT 282.120000 515.540000 283.320000 516.020000 ;
        RECT 282.120000 493.780000 283.320000 494.260000 ;
        RECT 282.120000 488.340000 283.320000 488.820000 ;
        RECT 282.120000 482.900000 283.320000 483.380000 ;
        RECT 282.120000 499.220000 283.320000 499.700000 ;
        RECT 282.120000 504.660000 283.320000 505.140000 ;
        RECT 282.120000 510.100000 283.320000 510.580000 ;
        RECT 327.120000 493.780000 328.320000 494.260000 ;
        RECT 327.120000 488.340000 328.320000 488.820000 ;
        RECT 327.120000 482.900000 328.320000 483.380000 ;
        RECT 327.120000 504.660000 328.320000 505.140000 ;
        RECT 327.120000 499.220000 328.320000 499.700000 ;
        RECT 327.120000 510.100000 328.320000 510.580000 ;
        RECT 282.120000 520.980000 283.320000 521.460000 ;
        RECT 282.120000 526.420000 283.320000 526.900000 ;
        RECT 282.120000 531.860000 283.320000 532.340000 ;
        RECT 282.120000 537.300000 283.320000 537.780000 ;
        RECT 327.120000 520.980000 328.320000 521.460000 ;
        RECT 327.120000 526.420000 328.320000 526.900000 ;
        RECT 327.120000 531.860000 328.320000 532.340000 ;
        RECT 327.120000 537.300000 328.320000 537.780000 ;
        RECT 372.120000 515.540000 373.320000 516.020000 ;
        RECT 372.120000 488.340000 373.320000 488.820000 ;
        RECT 372.120000 482.900000 373.320000 483.380000 ;
        RECT 372.120000 493.780000 373.320000 494.260000 ;
        RECT 372.120000 499.220000 373.320000 499.700000 ;
        RECT 372.120000 504.660000 373.320000 505.140000 ;
        RECT 372.120000 510.100000 373.320000 510.580000 ;
        RECT 372.120000 537.300000 373.320000 537.780000 ;
        RECT 372.120000 520.980000 373.320000 521.460000 ;
        RECT 372.120000 526.420000 373.320000 526.900000 ;
        RECT 372.120000 531.860000 373.320000 532.340000 ;
        RECT 417.120000 417.620000 418.320000 418.100000 ;
        RECT 417.120000 423.060000 418.320000 423.540000 ;
        RECT 417.120000 428.500000 418.320000 428.980000 ;
        RECT 417.120000 444.820000 418.320000 445.300000 ;
        RECT 417.120000 433.940000 418.320000 434.420000 ;
        RECT 417.120000 439.380000 418.320000 439.860000 ;
        RECT 462.120000 417.620000 463.320000 418.100000 ;
        RECT 462.120000 423.060000 463.320000 423.540000 ;
        RECT 462.120000 428.500000 463.320000 428.980000 ;
        RECT 462.120000 433.940000 463.320000 434.420000 ;
        RECT 462.120000 439.380000 463.320000 439.860000 ;
        RECT 462.120000 444.820000 463.320000 445.300000 ;
        RECT 417.120000 461.140000 418.320000 461.620000 ;
        RECT 417.120000 455.700000 418.320000 456.180000 ;
        RECT 417.120000 450.260000 418.320000 450.740000 ;
        RECT 417.120000 472.020000 418.320000 472.500000 ;
        RECT 417.120000 466.580000 418.320000 467.060000 ;
        RECT 417.120000 477.460000 418.320000 477.940000 ;
        RECT 462.120000 461.140000 463.320000 461.620000 ;
        RECT 462.120000 455.700000 463.320000 456.180000 ;
        RECT 462.120000 450.260000 463.320000 450.740000 ;
        RECT 462.120000 472.020000 463.320000 472.500000 ;
        RECT 462.120000 466.580000 463.320000 467.060000 ;
        RECT 462.120000 477.460000 463.320000 477.940000 ;
        RECT 507.120000 428.500000 508.320000 428.980000 ;
        RECT 507.120000 417.620000 508.320000 418.100000 ;
        RECT 507.120000 423.060000 508.320000 423.540000 ;
        RECT 507.120000 433.940000 508.320000 434.420000 ;
        RECT 507.120000 439.380000 508.320000 439.860000 ;
        RECT 507.120000 444.820000 508.320000 445.300000 ;
        RECT 543.400000 428.500000 544.600000 428.980000 ;
        RECT 543.400000 423.060000 544.600000 423.540000 ;
        RECT 543.400000 417.620000 544.600000 418.100000 ;
        RECT 543.400000 444.820000 544.600000 445.300000 ;
        RECT 543.400000 439.380000 544.600000 439.860000 ;
        RECT 543.400000 433.940000 544.600000 434.420000 ;
        RECT 507.120000 450.260000 508.320000 450.740000 ;
        RECT 507.120000 455.700000 508.320000 456.180000 ;
        RECT 507.120000 461.140000 508.320000 461.620000 ;
        RECT 507.120000 477.460000 508.320000 477.940000 ;
        RECT 507.120000 472.020000 508.320000 472.500000 ;
        RECT 507.120000 466.580000 508.320000 467.060000 ;
        RECT 543.400000 461.140000 544.600000 461.620000 ;
        RECT 543.400000 455.700000 544.600000 456.180000 ;
        RECT 543.400000 450.260000 544.600000 450.740000 ;
        RECT 543.400000 477.460000 544.600000 477.940000 ;
        RECT 543.400000 472.020000 544.600000 472.500000 ;
        RECT 543.400000 466.580000 544.600000 467.060000 ;
        RECT 462.120000 515.540000 463.320000 516.020000 ;
        RECT 417.120000 515.540000 418.320000 516.020000 ;
        RECT 417.120000 493.780000 418.320000 494.260000 ;
        RECT 417.120000 488.340000 418.320000 488.820000 ;
        RECT 417.120000 482.900000 418.320000 483.380000 ;
        RECT 417.120000 499.220000 418.320000 499.700000 ;
        RECT 417.120000 504.660000 418.320000 505.140000 ;
        RECT 417.120000 510.100000 418.320000 510.580000 ;
        RECT 462.120000 493.780000 463.320000 494.260000 ;
        RECT 462.120000 488.340000 463.320000 488.820000 ;
        RECT 462.120000 482.900000 463.320000 483.380000 ;
        RECT 462.120000 504.660000 463.320000 505.140000 ;
        RECT 462.120000 499.220000 463.320000 499.700000 ;
        RECT 462.120000 510.100000 463.320000 510.580000 ;
        RECT 417.120000 520.980000 418.320000 521.460000 ;
        RECT 417.120000 526.420000 418.320000 526.900000 ;
        RECT 417.120000 531.860000 418.320000 532.340000 ;
        RECT 417.120000 537.300000 418.320000 537.780000 ;
        RECT 462.120000 520.980000 463.320000 521.460000 ;
        RECT 462.120000 526.420000 463.320000 526.900000 ;
        RECT 462.120000 531.860000 463.320000 532.340000 ;
        RECT 462.120000 537.300000 463.320000 537.780000 ;
        RECT 543.400000 515.540000 544.600000 516.020000 ;
        RECT 507.120000 515.540000 508.320000 516.020000 ;
        RECT 507.120000 488.340000 508.320000 488.820000 ;
        RECT 507.120000 482.900000 508.320000 483.380000 ;
        RECT 507.120000 493.780000 508.320000 494.260000 ;
        RECT 507.120000 499.220000 508.320000 499.700000 ;
        RECT 507.120000 504.660000 508.320000 505.140000 ;
        RECT 507.120000 510.100000 508.320000 510.580000 ;
        RECT 543.400000 493.780000 544.600000 494.260000 ;
        RECT 543.400000 488.340000 544.600000 488.820000 ;
        RECT 543.400000 482.900000 544.600000 483.380000 ;
        RECT 543.400000 510.100000 544.600000 510.580000 ;
        RECT 543.400000 504.660000 544.600000 505.140000 ;
        RECT 543.400000 499.220000 544.600000 499.700000 ;
        RECT 507.120000 526.420000 508.320000 526.900000 ;
        RECT 507.120000 520.980000 508.320000 521.460000 ;
        RECT 507.120000 531.860000 508.320000 532.340000 ;
        RECT 507.120000 537.300000 508.320000 537.780000 ;
        RECT 543.400000 531.860000 544.600000 532.340000 ;
        RECT 543.400000 526.420000 544.600000 526.900000 ;
        RECT 543.400000 520.980000 544.600000 521.460000 ;
        RECT 543.400000 537.300000 544.600000 537.780000 ;
      LAYER met4 ;
        RECT 507.120000 5.430000 508.320000 543.160000 ;
        RECT 462.120000 5.430000 463.320000 543.160000 ;
        RECT 417.120000 5.430000 418.320000 543.160000 ;
        RECT 372.120000 5.430000 373.320000 543.160000 ;
        RECT 327.120000 5.430000 328.320000 543.160000 ;
        RECT 282.120000 5.430000 283.320000 543.160000 ;
        RECT 237.120000 5.430000 238.320000 543.160000 ;
        RECT 192.120000 5.430000 193.320000 543.160000 ;
        RECT 147.120000 5.430000 148.320000 543.160000 ;
        RECT 102.120000 5.430000 103.320000 543.160000 ;
        RECT 57.120000 5.430000 58.320000 543.160000 ;
        RECT 12.120000 5.430000 13.320000 543.160000 ;
        RECT 543.400000 0.000000 544.600000 549.780000 ;
        RECT 5.560000 0.000000 6.760000 549.780000 ;
    END
# end of P/G power stripe data as pin

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 548.960000 544.160000 550.160000 545.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 544.160000 1.200000 545.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 548.960000 3.230000 550.160000 4.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 3.230000 1.200000 4.430000 ;
    END
    PORT
      LAYER met4 ;
        RECT 545.600000 548.580000 546.800000 549.780000 ;
    END
    PORT
      LAYER met4 ;
        RECT 545.600000 0.000000 546.800000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 3.360000 548.580000 4.560000 549.780000 ;
    END
    PORT
      LAYER met4 ;
        RECT 3.360000 0.000000 4.560000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 3.230000 550.160000 4.430000 ;
        RECT 0.000000 544.160000 550.160000 545.360000 ;
        RECT 3.360000 34.100000 4.560000 34.580000 ;
        RECT 9.955000 34.100000 11.320000 34.580000 ;
        RECT 55.120000 34.100000 56.320000 34.580000 ;
        RECT 3.360000 12.340000 4.560000 12.820000 ;
        RECT 9.955000 12.340000 11.320000 12.820000 ;
        RECT 3.360000 23.220000 4.560000 23.700000 ;
        RECT 9.955000 23.220000 11.320000 23.700000 ;
        RECT 3.360000 17.780000 4.560000 18.260000 ;
        RECT 9.955000 17.780000 11.320000 18.260000 ;
        RECT 3.360000 28.660000 4.560000 29.140000 ;
        RECT 9.955000 28.660000 11.320000 29.140000 ;
        RECT 55.120000 28.660000 56.320000 29.140000 ;
        RECT 55.120000 23.220000 56.320000 23.700000 ;
        RECT 55.120000 17.780000 56.320000 18.260000 ;
        RECT 55.120000 12.340000 56.320000 12.820000 ;
        RECT 3.360000 39.540000 4.560000 40.020000 ;
        RECT 9.955000 39.540000 11.320000 40.020000 ;
        RECT 3.360000 50.420000 4.560000 50.900000 ;
        RECT 9.955000 50.420000 11.320000 50.900000 ;
        RECT 3.360000 44.980000 4.560000 45.460000 ;
        RECT 9.955000 44.980000 11.320000 45.460000 ;
        RECT 3.360000 55.860000 4.560000 56.340000 ;
        RECT 9.955000 55.860000 11.320000 56.340000 ;
        RECT 3.360000 66.740000 4.560000 67.220000 ;
        RECT 9.955000 66.740000 11.320000 67.220000 ;
        RECT 3.360000 61.300000 4.560000 61.780000 ;
        RECT 9.955000 61.300000 11.320000 61.780000 ;
        RECT 55.120000 39.540000 56.320000 40.020000 ;
        RECT 55.120000 44.980000 56.320000 45.460000 ;
        RECT 55.120000 50.420000 56.320000 50.900000 ;
        RECT 55.120000 66.740000 56.320000 67.220000 ;
        RECT 55.120000 61.300000 56.320000 61.780000 ;
        RECT 55.120000 55.860000 56.320000 56.340000 ;
        RECT 100.120000 34.100000 101.320000 34.580000 ;
        RECT 100.120000 28.660000 101.320000 29.140000 ;
        RECT 100.120000 23.220000 101.320000 23.700000 ;
        RECT 100.120000 17.780000 101.320000 18.260000 ;
        RECT 100.120000 12.340000 101.320000 12.820000 ;
        RECT 100.120000 66.740000 101.320000 67.220000 ;
        RECT 100.120000 61.300000 101.320000 61.780000 ;
        RECT 100.120000 39.540000 101.320000 40.020000 ;
        RECT 100.120000 44.980000 101.320000 45.460000 ;
        RECT 100.120000 50.420000 101.320000 50.900000 ;
        RECT 100.120000 55.860000 101.320000 56.340000 ;
        RECT 3.360000 72.180000 4.560000 72.660000 ;
        RECT 9.955000 72.180000 11.320000 72.660000 ;
        RECT 3.360000 83.060000 4.560000 83.540000 ;
        RECT 9.955000 83.060000 11.320000 83.540000 ;
        RECT 3.360000 77.620000 4.560000 78.100000 ;
        RECT 9.955000 77.620000 11.320000 78.100000 ;
        RECT 3.360000 93.940000 4.560000 94.420000 ;
        RECT 9.955000 93.940000 11.320000 94.420000 ;
        RECT 3.360000 88.500000 4.560000 88.980000 ;
        RECT 9.955000 88.500000 11.320000 88.980000 ;
        RECT 3.360000 99.380000 4.560000 99.860000 ;
        RECT 9.955000 99.380000 11.320000 99.860000 ;
        RECT 55.120000 72.180000 56.320000 72.660000 ;
        RECT 55.120000 77.620000 56.320000 78.100000 ;
        RECT 55.120000 83.060000 56.320000 83.540000 ;
        RECT 55.120000 99.380000 56.320000 99.860000 ;
        RECT 55.120000 93.940000 56.320000 94.420000 ;
        RECT 55.120000 88.500000 56.320000 88.980000 ;
        RECT 3.360000 110.260000 4.560000 110.740000 ;
        RECT 9.955000 110.260000 11.320000 110.740000 ;
        RECT 3.360000 104.820000 4.560000 105.300000 ;
        RECT 9.955000 104.820000 11.320000 105.300000 ;
        RECT 3.360000 115.700000 4.560000 116.180000 ;
        RECT 9.955000 115.700000 11.320000 116.180000 ;
        RECT 3.360000 126.580000 4.560000 127.060000 ;
        RECT 9.955000 126.580000 11.320000 127.060000 ;
        RECT 3.360000 121.140000 4.560000 121.620000 ;
        RECT 9.955000 121.140000 11.320000 121.620000 ;
        RECT 3.360000 132.020000 4.560000 132.500000 ;
        RECT 9.955000 132.020000 11.320000 132.500000 ;
        RECT 55.120000 104.820000 56.320000 105.300000 ;
        RECT 55.120000 110.260000 56.320000 110.740000 ;
        RECT 55.120000 115.700000 56.320000 116.180000 ;
        RECT 55.120000 132.020000 56.320000 132.500000 ;
        RECT 55.120000 126.580000 56.320000 127.060000 ;
        RECT 55.120000 121.140000 56.320000 121.620000 ;
        RECT 100.120000 99.380000 101.320000 99.860000 ;
        RECT 100.120000 93.940000 101.320000 94.420000 ;
        RECT 100.120000 88.500000 101.320000 88.980000 ;
        RECT 100.120000 72.180000 101.320000 72.660000 ;
        RECT 100.120000 77.620000 101.320000 78.100000 ;
        RECT 100.120000 83.060000 101.320000 83.540000 ;
        RECT 100.120000 132.020000 101.320000 132.500000 ;
        RECT 100.120000 126.580000 101.320000 127.060000 ;
        RECT 100.120000 104.820000 101.320000 105.300000 ;
        RECT 100.120000 110.260000 101.320000 110.740000 ;
        RECT 100.120000 115.700000 101.320000 116.180000 ;
        RECT 100.120000 121.140000 101.320000 121.620000 ;
        RECT 190.120000 34.100000 191.320000 34.580000 ;
        RECT 145.120000 34.100000 146.320000 34.580000 ;
        RECT 145.120000 28.660000 146.320000 29.140000 ;
        RECT 145.120000 23.220000 146.320000 23.700000 ;
        RECT 145.120000 17.780000 146.320000 18.260000 ;
        RECT 145.120000 12.340000 146.320000 12.820000 ;
        RECT 190.120000 28.660000 191.320000 29.140000 ;
        RECT 190.120000 23.220000 191.320000 23.700000 ;
        RECT 190.120000 17.780000 191.320000 18.260000 ;
        RECT 190.120000 12.340000 191.320000 12.820000 ;
        RECT 145.120000 39.540000 146.320000 40.020000 ;
        RECT 145.120000 44.980000 146.320000 45.460000 ;
        RECT 145.120000 50.420000 146.320000 50.900000 ;
        RECT 145.120000 66.740000 146.320000 67.220000 ;
        RECT 145.120000 61.300000 146.320000 61.780000 ;
        RECT 145.120000 55.860000 146.320000 56.340000 ;
        RECT 190.120000 39.540000 191.320000 40.020000 ;
        RECT 190.120000 44.980000 191.320000 45.460000 ;
        RECT 190.120000 50.420000 191.320000 50.900000 ;
        RECT 190.120000 66.740000 191.320000 67.220000 ;
        RECT 190.120000 61.300000 191.320000 61.780000 ;
        RECT 190.120000 55.860000 191.320000 56.340000 ;
        RECT 235.120000 34.100000 236.320000 34.580000 ;
        RECT 235.120000 28.660000 236.320000 29.140000 ;
        RECT 235.120000 23.220000 236.320000 23.700000 ;
        RECT 235.120000 17.780000 236.320000 18.260000 ;
        RECT 235.120000 12.340000 236.320000 12.820000 ;
        RECT 235.120000 50.420000 236.320000 50.900000 ;
        RECT 235.120000 44.980000 236.320000 45.460000 ;
        RECT 235.120000 39.540000 236.320000 40.020000 ;
        RECT 235.120000 66.740000 236.320000 67.220000 ;
        RECT 235.120000 55.860000 236.320000 56.340000 ;
        RECT 235.120000 61.300000 236.320000 61.780000 ;
        RECT 145.120000 72.180000 146.320000 72.660000 ;
        RECT 145.120000 77.620000 146.320000 78.100000 ;
        RECT 145.120000 83.060000 146.320000 83.540000 ;
        RECT 145.120000 99.380000 146.320000 99.860000 ;
        RECT 145.120000 93.940000 146.320000 94.420000 ;
        RECT 145.120000 88.500000 146.320000 88.980000 ;
        RECT 190.120000 72.180000 191.320000 72.660000 ;
        RECT 190.120000 77.620000 191.320000 78.100000 ;
        RECT 190.120000 83.060000 191.320000 83.540000 ;
        RECT 190.120000 99.380000 191.320000 99.860000 ;
        RECT 190.120000 93.940000 191.320000 94.420000 ;
        RECT 190.120000 88.500000 191.320000 88.980000 ;
        RECT 145.120000 104.820000 146.320000 105.300000 ;
        RECT 145.120000 110.260000 146.320000 110.740000 ;
        RECT 145.120000 115.700000 146.320000 116.180000 ;
        RECT 145.120000 132.020000 146.320000 132.500000 ;
        RECT 145.120000 126.580000 146.320000 127.060000 ;
        RECT 145.120000 121.140000 146.320000 121.620000 ;
        RECT 190.120000 104.820000 191.320000 105.300000 ;
        RECT 190.120000 110.260000 191.320000 110.740000 ;
        RECT 190.120000 115.700000 191.320000 116.180000 ;
        RECT 190.120000 132.020000 191.320000 132.500000 ;
        RECT 190.120000 126.580000 191.320000 127.060000 ;
        RECT 190.120000 121.140000 191.320000 121.620000 ;
        RECT 235.120000 83.060000 236.320000 83.540000 ;
        RECT 235.120000 77.620000 236.320000 78.100000 ;
        RECT 235.120000 72.180000 236.320000 72.660000 ;
        RECT 235.120000 99.380000 236.320000 99.860000 ;
        RECT 235.120000 93.940000 236.320000 94.420000 ;
        RECT 235.120000 88.500000 236.320000 88.980000 ;
        RECT 235.120000 115.700000 236.320000 116.180000 ;
        RECT 235.120000 110.260000 236.320000 110.740000 ;
        RECT 235.120000 104.820000 236.320000 105.300000 ;
        RECT 235.120000 132.020000 236.320000 132.500000 ;
        RECT 235.120000 121.140000 236.320000 121.620000 ;
        RECT 235.120000 126.580000 236.320000 127.060000 ;
        RECT 3.360000 142.900000 4.560000 143.380000 ;
        RECT 9.955000 142.900000 11.320000 143.380000 ;
        RECT 3.360000 137.460000 4.560000 137.940000 ;
        RECT 9.955000 137.460000 11.320000 137.940000 ;
        RECT 3.360000 153.780000 4.560000 154.260000 ;
        RECT 9.955000 153.780000 11.320000 154.260000 ;
        RECT 3.360000 148.340000 4.560000 148.820000 ;
        RECT 9.955000 148.340000 11.320000 148.820000 ;
        RECT 3.360000 159.220000 4.560000 159.700000 ;
        RECT 9.955000 159.220000 11.320000 159.700000 ;
        RECT 3.360000 170.100000 4.560000 170.580000 ;
        RECT 9.955000 170.100000 11.320000 170.580000 ;
        RECT 3.360000 164.660000 4.560000 165.140000 ;
        RECT 9.955000 164.660000 11.320000 165.140000 ;
        RECT 55.120000 137.460000 56.320000 137.940000 ;
        RECT 55.120000 142.900000 56.320000 143.380000 ;
        RECT 55.120000 148.340000 56.320000 148.820000 ;
        RECT 55.120000 153.780000 56.320000 154.260000 ;
        RECT 55.120000 170.100000 56.320000 170.580000 ;
        RECT 55.120000 164.660000 56.320000 165.140000 ;
        RECT 55.120000 159.220000 56.320000 159.700000 ;
        RECT 3.360000 175.540000 4.560000 176.020000 ;
        RECT 9.955000 175.540000 11.320000 176.020000 ;
        RECT 3.360000 186.420000 4.560000 186.900000 ;
        RECT 9.955000 186.420000 11.320000 186.900000 ;
        RECT 3.360000 180.980000 4.560000 181.460000 ;
        RECT 9.955000 180.980000 11.320000 181.460000 ;
        RECT 3.360000 197.300000 4.560000 197.780000 ;
        RECT 9.955000 197.300000 11.320000 197.780000 ;
        RECT 3.360000 191.860000 4.560000 192.340000 ;
        RECT 9.955000 191.860000 11.320000 192.340000 ;
        RECT 3.360000 202.740000 4.560000 203.220000 ;
        RECT 9.955000 202.740000 11.320000 203.220000 ;
        RECT 55.120000 175.540000 56.320000 176.020000 ;
        RECT 55.120000 180.980000 56.320000 181.460000 ;
        RECT 55.120000 186.420000 56.320000 186.900000 ;
        RECT 55.120000 202.740000 56.320000 203.220000 ;
        RECT 55.120000 197.300000 56.320000 197.780000 ;
        RECT 55.120000 191.860000 56.320000 192.340000 ;
        RECT 100.120000 170.100000 101.320000 170.580000 ;
        RECT 100.120000 164.660000 101.320000 165.140000 ;
        RECT 100.120000 159.220000 101.320000 159.700000 ;
        RECT 100.120000 137.460000 101.320000 137.940000 ;
        RECT 100.120000 142.900000 101.320000 143.380000 ;
        RECT 100.120000 148.340000 101.320000 148.820000 ;
        RECT 100.120000 153.780000 101.320000 154.260000 ;
        RECT 100.120000 202.740000 101.320000 203.220000 ;
        RECT 100.120000 197.300000 101.320000 197.780000 ;
        RECT 100.120000 191.860000 101.320000 192.340000 ;
        RECT 100.120000 175.540000 101.320000 176.020000 ;
        RECT 100.120000 180.980000 101.320000 181.460000 ;
        RECT 100.120000 186.420000 101.320000 186.900000 ;
        RECT 3.360000 213.620000 4.560000 214.100000 ;
        RECT 9.955000 213.620000 11.320000 214.100000 ;
        RECT 3.360000 208.180000 4.560000 208.660000 ;
        RECT 9.955000 208.180000 11.320000 208.660000 ;
        RECT 3.360000 219.060000 4.560000 219.540000 ;
        RECT 9.955000 219.060000 11.320000 219.540000 ;
        RECT 3.360000 229.940000 4.560000 230.420000 ;
        RECT 9.955000 229.940000 11.320000 230.420000 ;
        RECT 3.360000 224.500000 4.560000 224.980000 ;
        RECT 9.955000 224.500000 11.320000 224.980000 ;
        RECT 3.360000 235.380000 4.560000 235.860000 ;
        RECT 9.955000 235.380000 11.320000 235.860000 ;
        RECT 55.120000 208.180000 56.320000 208.660000 ;
        RECT 55.120000 213.620000 56.320000 214.100000 ;
        RECT 55.120000 219.060000 56.320000 219.540000 ;
        RECT 55.120000 235.380000 56.320000 235.860000 ;
        RECT 55.120000 229.940000 56.320000 230.420000 ;
        RECT 55.120000 224.500000 56.320000 224.980000 ;
        RECT 3.360000 246.260000 4.560000 246.740000 ;
        RECT 9.955000 246.260000 11.320000 246.740000 ;
        RECT 3.360000 240.820000 4.560000 241.300000 ;
        RECT 9.955000 240.820000 11.320000 241.300000 ;
        RECT 3.360000 257.140000 4.560000 257.620000 ;
        RECT 9.955000 257.140000 11.320000 257.620000 ;
        RECT 3.360000 251.700000 4.560000 252.180000 ;
        RECT 9.955000 251.700000 11.320000 252.180000 ;
        RECT 3.360000 262.580000 4.560000 263.060000 ;
        RECT 9.955000 262.580000 11.320000 263.060000 ;
        RECT 3.360000 273.460000 4.560000 273.940000 ;
        RECT 9.955000 273.460000 11.320000 273.940000 ;
        RECT 3.360000 268.020000 4.560000 268.500000 ;
        RECT 9.955000 268.020000 11.320000 268.500000 ;
        RECT 55.120000 240.820000 56.320000 241.300000 ;
        RECT 55.120000 246.260000 56.320000 246.740000 ;
        RECT 55.120000 251.700000 56.320000 252.180000 ;
        RECT 55.120000 257.140000 56.320000 257.620000 ;
        RECT 55.120000 273.460000 56.320000 273.940000 ;
        RECT 55.120000 268.020000 56.320000 268.500000 ;
        RECT 55.120000 262.580000 56.320000 263.060000 ;
        RECT 100.120000 235.380000 101.320000 235.860000 ;
        RECT 100.120000 229.940000 101.320000 230.420000 ;
        RECT 100.120000 208.180000 101.320000 208.660000 ;
        RECT 100.120000 213.620000 101.320000 214.100000 ;
        RECT 100.120000 219.060000 101.320000 219.540000 ;
        RECT 100.120000 224.500000 101.320000 224.980000 ;
        RECT 100.120000 273.460000 101.320000 273.940000 ;
        RECT 100.120000 268.020000 101.320000 268.500000 ;
        RECT 100.120000 262.580000 101.320000 263.060000 ;
        RECT 100.120000 240.820000 101.320000 241.300000 ;
        RECT 100.120000 246.260000 101.320000 246.740000 ;
        RECT 100.120000 251.700000 101.320000 252.180000 ;
        RECT 100.120000 257.140000 101.320000 257.620000 ;
        RECT 145.120000 137.460000 146.320000 137.940000 ;
        RECT 145.120000 142.900000 146.320000 143.380000 ;
        RECT 145.120000 148.340000 146.320000 148.820000 ;
        RECT 145.120000 153.780000 146.320000 154.260000 ;
        RECT 145.120000 170.100000 146.320000 170.580000 ;
        RECT 145.120000 164.660000 146.320000 165.140000 ;
        RECT 145.120000 159.220000 146.320000 159.700000 ;
        RECT 190.120000 137.460000 191.320000 137.940000 ;
        RECT 190.120000 142.900000 191.320000 143.380000 ;
        RECT 190.120000 148.340000 191.320000 148.820000 ;
        RECT 190.120000 153.780000 191.320000 154.260000 ;
        RECT 190.120000 170.100000 191.320000 170.580000 ;
        RECT 190.120000 164.660000 191.320000 165.140000 ;
        RECT 190.120000 159.220000 191.320000 159.700000 ;
        RECT 145.120000 175.540000 146.320000 176.020000 ;
        RECT 145.120000 180.980000 146.320000 181.460000 ;
        RECT 145.120000 186.420000 146.320000 186.900000 ;
        RECT 145.120000 202.740000 146.320000 203.220000 ;
        RECT 145.120000 197.300000 146.320000 197.780000 ;
        RECT 145.120000 191.860000 146.320000 192.340000 ;
        RECT 190.120000 175.540000 191.320000 176.020000 ;
        RECT 190.120000 180.980000 191.320000 181.460000 ;
        RECT 190.120000 186.420000 191.320000 186.900000 ;
        RECT 190.120000 202.740000 191.320000 203.220000 ;
        RECT 190.120000 197.300000 191.320000 197.780000 ;
        RECT 190.120000 191.860000 191.320000 192.340000 ;
        RECT 235.120000 153.780000 236.320000 154.260000 ;
        RECT 235.120000 148.340000 236.320000 148.820000 ;
        RECT 235.120000 142.900000 236.320000 143.380000 ;
        RECT 235.120000 137.460000 236.320000 137.940000 ;
        RECT 235.120000 170.100000 236.320000 170.580000 ;
        RECT 235.120000 164.660000 236.320000 165.140000 ;
        RECT 235.120000 159.220000 236.320000 159.700000 ;
        RECT 235.120000 186.420000 236.320000 186.900000 ;
        RECT 235.120000 180.980000 236.320000 181.460000 ;
        RECT 235.120000 175.540000 236.320000 176.020000 ;
        RECT 235.120000 202.740000 236.320000 203.220000 ;
        RECT 235.120000 197.300000 236.320000 197.780000 ;
        RECT 235.120000 191.860000 236.320000 192.340000 ;
        RECT 145.120000 208.180000 146.320000 208.660000 ;
        RECT 145.120000 213.620000 146.320000 214.100000 ;
        RECT 145.120000 219.060000 146.320000 219.540000 ;
        RECT 145.120000 235.380000 146.320000 235.860000 ;
        RECT 145.120000 229.940000 146.320000 230.420000 ;
        RECT 145.120000 224.500000 146.320000 224.980000 ;
        RECT 190.120000 208.180000 191.320000 208.660000 ;
        RECT 190.120000 213.620000 191.320000 214.100000 ;
        RECT 190.120000 219.060000 191.320000 219.540000 ;
        RECT 190.120000 235.380000 191.320000 235.860000 ;
        RECT 190.120000 229.940000 191.320000 230.420000 ;
        RECT 190.120000 224.500000 191.320000 224.980000 ;
        RECT 145.120000 240.820000 146.320000 241.300000 ;
        RECT 145.120000 246.260000 146.320000 246.740000 ;
        RECT 145.120000 251.700000 146.320000 252.180000 ;
        RECT 145.120000 257.140000 146.320000 257.620000 ;
        RECT 145.120000 273.460000 146.320000 273.940000 ;
        RECT 145.120000 268.020000 146.320000 268.500000 ;
        RECT 145.120000 262.580000 146.320000 263.060000 ;
        RECT 190.120000 240.820000 191.320000 241.300000 ;
        RECT 190.120000 246.260000 191.320000 246.740000 ;
        RECT 190.120000 251.700000 191.320000 252.180000 ;
        RECT 190.120000 257.140000 191.320000 257.620000 ;
        RECT 190.120000 273.460000 191.320000 273.940000 ;
        RECT 190.120000 268.020000 191.320000 268.500000 ;
        RECT 190.120000 262.580000 191.320000 263.060000 ;
        RECT 235.120000 219.060000 236.320000 219.540000 ;
        RECT 235.120000 213.620000 236.320000 214.100000 ;
        RECT 235.120000 208.180000 236.320000 208.660000 ;
        RECT 235.120000 235.380000 236.320000 235.860000 ;
        RECT 235.120000 224.500000 236.320000 224.980000 ;
        RECT 235.120000 229.940000 236.320000 230.420000 ;
        RECT 235.120000 257.140000 236.320000 257.620000 ;
        RECT 235.120000 251.700000 236.320000 252.180000 ;
        RECT 235.120000 246.260000 236.320000 246.740000 ;
        RECT 235.120000 240.820000 236.320000 241.300000 ;
        RECT 235.120000 273.460000 236.320000 273.940000 ;
        RECT 235.120000 268.020000 236.320000 268.500000 ;
        RECT 235.120000 262.580000 236.320000 263.060000 ;
        RECT 325.120000 34.100000 326.320000 34.580000 ;
        RECT 280.120000 34.100000 281.320000 34.580000 ;
        RECT 280.120000 28.660000 281.320000 29.140000 ;
        RECT 280.120000 23.220000 281.320000 23.700000 ;
        RECT 280.120000 17.780000 281.320000 18.260000 ;
        RECT 280.120000 12.340000 281.320000 12.820000 ;
        RECT 325.120000 28.660000 326.320000 29.140000 ;
        RECT 325.120000 23.220000 326.320000 23.700000 ;
        RECT 325.120000 17.780000 326.320000 18.260000 ;
        RECT 325.120000 12.340000 326.320000 12.820000 ;
        RECT 280.120000 39.540000 281.320000 40.020000 ;
        RECT 280.120000 44.980000 281.320000 45.460000 ;
        RECT 280.120000 50.420000 281.320000 50.900000 ;
        RECT 280.120000 66.740000 281.320000 67.220000 ;
        RECT 280.120000 61.300000 281.320000 61.780000 ;
        RECT 280.120000 55.860000 281.320000 56.340000 ;
        RECT 325.120000 39.540000 326.320000 40.020000 ;
        RECT 325.120000 44.980000 326.320000 45.460000 ;
        RECT 325.120000 50.420000 326.320000 50.900000 ;
        RECT 325.120000 66.740000 326.320000 67.220000 ;
        RECT 325.120000 61.300000 326.320000 61.780000 ;
        RECT 325.120000 55.860000 326.320000 56.340000 ;
        RECT 370.120000 34.100000 371.320000 34.580000 ;
        RECT 370.120000 28.660000 371.320000 29.140000 ;
        RECT 370.120000 23.220000 371.320000 23.700000 ;
        RECT 370.120000 17.780000 371.320000 18.260000 ;
        RECT 370.120000 12.340000 371.320000 12.820000 ;
        RECT 370.120000 50.420000 371.320000 50.900000 ;
        RECT 370.120000 44.980000 371.320000 45.460000 ;
        RECT 370.120000 39.540000 371.320000 40.020000 ;
        RECT 370.120000 66.740000 371.320000 67.220000 ;
        RECT 370.120000 55.860000 371.320000 56.340000 ;
        RECT 370.120000 61.300000 371.320000 61.780000 ;
        RECT 280.120000 72.180000 281.320000 72.660000 ;
        RECT 280.120000 77.620000 281.320000 78.100000 ;
        RECT 280.120000 83.060000 281.320000 83.540000 ;
        RECT 280.120000 99.380000 281.320000 99.860000 ;
        RECT 280.120000 93.940000 281.320000 94.420000 ;
        RECT 280.120000 88.500000 281.320000 88.980000 ;
        RECT 325.120000 72.180000 326.320000 72.660000 ;
        RECT 325.120000 77.620000 326.320000 78.100000 ;
        RECT 325.120000 83.060000 326.320000 83.540000 ;
        RECT 325.120000 99.380000 326.320000 99.860000 ;
        RECT 325.120000 93.940000 326.320000 94.420000 ;
        RECT 325.120000 88.500000 326.320000 88.980000 ;
        RECT 280.120000 104.820000 281.320000 105.300000 ;
        RECT 280.120000 110.260000 281.320000 110.740000 ;
        RECT 280.120000 115.700000 281.320000 116.180000 ;
        RECT 280.120000 132.020000 281.320000 132.500000 ;
        RECT 280.120000 126.580000 281.320000 127.060000 ;
        RECT 280.120000 121.140000 281.320000 121.620000 ;
        RECT 325.120000 104.820000 326.320000 105.300000 ;
        RECT 325.120000 110.260000 326.320000 110.740000 ;
        RECT 325.120000 115.700000 326.320000 116.180000 ;
        RECT 325.120000 132.020000 326.320000 132.500000 ;
        RECT 325.120000 126.580000 326.320000 127.060000 ;
        RECT 325.120000 121.140000 326.320000 121.620000 ;
        RECT 370.120000 83.060000 371.320000 83.540000 ;
        RECT 370.120000 77.620000 371.320000 78.100000 ;
        RECT 370.120000 72.180000 371.320000 72.660000 ;
        RECT 370.120000 99.380000 371.320000 99.860000 ;
        RECT 370.120000 93.940000 371.320000 94.420000 ;
        RECT 370.120000 88.500000 371.320000 88.980000 ;
        RECT 370.120000 115.700000 371.320000 116.180000 ;
        RECT 370.120000 110.260000 371.320000 110.740000 ;
        RECT 370.120000 104.820000 371.320000 105.300000 ;
        RECT 370.120000 132.020000 371.320000 132.500000 ;
        RECT 370.120000 121.140000 371.320000 121.620000 ;
        RECT 370.120000 126.580000 371.320000 127.060000 ;
        RECT 460.120000 34.100000 461.320000 34.580000 ;
        RECT 415.120000 34.100000 416.320000 34.580000 ;
        RECT 415.120000 28.660000 416.320000 29.140000 ;
        RECT 415.120000 23.220000 416.320000 23.700000 ;
        RECT 415.120000 17.780000 416.320000 18.260000 ;
        RECT 415.120000 12.340000 416.320000 12.820000 ;
        RECT 460.120000 28.660000 461.320000 29.140000 ;
        RECT 460.120000 23.220000 461.320000 23.700000 ;
        RECT 460.120000 17.780000 461.320000 18.260000 ;
        RECT 460.120000 12.340000 461.320000 12.820000 ;
        RECT 415.120000 39.540000 416.320000 40.020000 ;
        RECT 415.120000 44.980000 416.320000 45.460000 ;
        RECT 415.120000 50.420000 416.320000 50.900000 ;
        RECT 415.120000 66.740000 416.320000 67.220000 ;
        RECT 415.120000 61.300000 416.320000 61.780000 ;
        RECT 415.120000 55.860000 416.320000 56.340000 ;
        RECT 460.120000 39.540000 461.320000 40.020000 ;
        RECT 460.120000 44.980000 461.320000 45.460000 ;
        RECT 460.120000 50.420000 461.320000 50.900000 ;
        RECT 460.120000 66.740000 461.320000 67.220000 ;
        RECT 460.120000 61.300000 461.320000 61.780000 ;
        RECT 460.120000 55.860000 461.320000 56.340000 ;
        RECT 545.600000 34.100000 546.800000 34.580000 ;
        RECT 505.120000 34.100000 506.320000 34.580000 ;
        RECT 505.120000 12.340000 506.320000 12.820000 ;
        RECT 505.120000 17.780000 506.320000 18.260000 ;
        RECT 505.120000 23.220000 506.320000 23.700000 ;
        RECT 505.120000 28.660000 506.320000 29.140000 ;
        RECT 545.600000 12.340000 546.800000 12.820000 ;
        RECT 545.600000 28.660000 546.800000 29.140000 ;
        RECT 545.600000 23.220000 546.800000 23.700000 ;
        RECT 545.600000 17.780000 546.800000 18.260000 ;
        RECT 505.120000 50.420000 506.320000 50.900000 ;
        RECT 505.120000 44.980000 506.320000 45.460000 ;
        RECT 505.120000 39.540000 506.320000 40.020000 ;
        RECT 505.120000 66.740000 506.320000 67.220000 ;
        RECT 505.120000 55.860000 506.320000 56.340000 ;
        RECT 505.120000 61.300000 506.320000 61.780000 ;
        RECT 545.600000 50.420000 546.800000 50.900000 ;
        RECT 545.600000 39.540000 546.800000 40.020000 ;
        RECT 545.600000 44.980000 546.800000 45.460000 ;
        RECT 545.600000 66.740000 546.800000 67.220000 ;
        RECT 545.600000 61.300000 546.800000 61.780000 ;
        RECT 545.600000 55.860000 546.800000 56.340000 ;
        RECT 415.120000 72.180000 416.320000 72.660000 ;
        RECT 415.120000 77.620000 416.320000 78.100000 ;
        RECT 415.120000 83.060000 416.320000 83.540000 ;
        RECT 415.120000 99.380000 416.320000 99.860000 ;
        RECT 415.120000 93.940000 416.320000 94.420000 ;
        RECT 415.120000 88.500000 416.320000 88.980000 ;
        RECT 460.120000 72.180000 461.320000 72.660000 ;
        RECT 460.120000 77.620000 461.320000 78.100000 ;
        RECT 460.120000 83.060000 461.320000 83.540000 ;
        RECT 460.120000 99.380000 461.320000 99.860000 ;
        RECT 460.120000 93.940000 461.320000 94.420000 ;
        RECT 460.120000 88.500000 461.320000 88.980000 ;
        RECT 415.120000 104.820000 416.320000 105.300000 ;
        RECT 415.120000 110.260000 416.320000 110.740000 ;
        RECT 415.120000 115.700000 416.320000 116.180000 ;
        RECT 415.120000 132.020000 416.320000 132.500000 ;
        RECT 415.120000 126.580000 416.320000 127.060000 ;
        RECT 415.120000 121.140000 416.320000 121.620000 ;
        RECT 460.120000 104.820000 461.320000 105.300000 ;
        RECT 460.120000 110.260000 461.320000 110.740000 ;
        RECT 460.120000 115.700000 461.320000 116.180000 ;
        RECT 460.120000 132.020000 461.320000 132.500000 ;
        RECT 460.120000 126.580000 461.320000 127.060000 ;
        RECT 460.120000 121.140000 461.320000 121.620000 ;
        RECT 505.120000 83.060000 506.320000 83.540000 ;
        RECT 505.120000 77.620000 506.320000 78.100000 ;
        RECT 505.120000 72.180000 506.320000 72.660000 ;
        RECT 505.120000 99.380000 506.320000 99.860000 ;
        RECT 505.120000 93.940000 506.320000 94.420000 ;
        RECT 505.120000 88.500000 506.320000 88.980000 ;
        RECT 545.600000 83.060000 546.800000 83.540000 ;
        RECT 545.600000 77.620000 546.800000 78.100000 ;
        RECT 545.600000 72.180000 546.800000 72.660000 ;
        RECT 545.600000 99.380000 546.800000 99.860000 ;
        RECT 545.600000 93.940000 546.800000 94.420000 ;
        RECT 545.600000 88.500000 546.800000 88.980000 ;
        RECT 505.120000 115.700000 506.320000 116.180000 ;
        RECT 505.120000 110.260000 506.320000 110.740000 ;
        RECT 505.120000 104.820000 506.320000 105.300000 ;
        RECT 505.120000 132.020000 506.320000 132.500000 ;
        RECT 505.120000 121.140000 506.320000 121.620000 ;
        RECT 505.120000 126.580000 506.320000 127.060000 ;
        RECT 545.600000 115.700000 546.800000 116.180000 ;
        RECT 545.600000 104.820000 546.800000 105.300000 ;
        RECT 545.600000 110.260000 546.800000 110.740000 ;
        RECT 545.600000 132.020000 546.800000 132.500000 ;
        RECT 545.600000 126.580000 546.800000 127.060000 ;
        RECT 545.600000 121.140000 546.800000 121.620000 ;
        RECT 280.120000 137.460000 281.320000 137.940000 ;
        RECT 280.120000 142.900000 281.320000 143.380000 ;
        RECT 280.120000 148.340000 281.320000 148.820000 ;
        RECT 280.120000 153.780000 281.320000 154.260000 ;
        RECT 280.120000 170.100000 281.320000 170.580000 ;
        RECT 280.120000 164.660000 281.320000 165.140000 ;
        RECT 280.120000 159.220000 281.320000 159.700000 ;
        RECT 325.120000 137.460000 326.320000 137.940000 ;
        RECT 325.120000 142.900000 326.320000 143.380000 ;
        RECT 325.120000 148.340000 326.320000 148.820000 ;
        RECT 325.120000 153.780000 326.320000 154.260000 ;
        RECT 325.120000 170.100000 326.320000 170.580000 ;
        RECT 325.120000 164.660000 326.320000 165.140000 ;
        RECT 325.120000 159.220000 326.320000 159.700000 ;
        RECT 280.120000 175.540000 281.320000 176.020000 ;
        RECT 280.120000 180.980000 281.320000 181.460000 ;
        RECT 280.120000 186.420000 281.320000 186.900000 ;
        RECT 280.120000 202.740000 281.320000 203.220000 ;
        RECT 280.120000 197.300000 281.320000 197.780000 ;
        RECT 280.120000 191.860000 281.320000 192.340000 ;
        RECT 325.120000 175.540000 326.320000 176.020000 ;
        RECT 325.120000 180.980000 326.320000 181.460000 ;
        RECT 325.120000 186.420000 326.320000 186.900000 ;
        RECT 325.120000 202.740000 326.320000 203.220000 ;
        RECT 325.120000 197.300000 326.320000 197.780000 ;
        RECT 325.120000 191.860000 326.320000 192.340000 ;
        RECT 370.120000 153.780000 371.320000 154.260000 ;
        RECT 370.120000 148.340000 371.320000 148.820000 ;
        RECT 370.120000 142.900000 371.320000 143.380000 ;
        RECT 370.120000 137.460000 371.320000 137.940000 ;
        RECT 370.120000 170.100000 371.320000 170.580000 ;
        RECT 370.120000 164.660000 371.320000 165.140000 ;
        RECT 370.120000 159.220000 371.320000 159.700000 ;
        RECT 370.120000 186.420000 371.320000 186.900000 ;
        RECT 370.120000 180.980000 371.320000 181.460000 ;
        RECT 370.120000 175.540000 371.320000 176.020000 ;
        RECT 370.120000 202.740000 371.320000 203.220000 ;
        RECT 370.120000 197.300000 371.320000 197.780000 ;
        RECT 370.120000 191.860000 371.320000 192.340000 ;
        RECT 280.120000 208.180000 281.320000 208.660000 ;
        RECT 280.120000 213.620000 281.320000 214.100000 ;
        RECT 280.120000 219.060000 281.320000 219.540000 ;
        RECT 280.120000 235.380000 281.320000 235.860000 ;
        RECT 280.120000 229.940000 281.320000 230.420000 ;
        RECT 280.120000 224.500000 281.320000 224.980000 ;
        RECT 325.120000 208.180000 326.320000 208.660000 ;
        RECT 325.120000 213.620000 326.320000 214.100000 ;
        RECT 325.120000 219.060000 326.320000 219.540000 ;
        RECT 325.120000 235.380000 326.320000 235.860000 ;
        RECT 325.120000 229.940000 326.320000 230.420000 ;
        RECT 325.120000 224.500000 326.320000 224.980000 ;
        RECT 280.120000 240.820000 281.320000 241.300000 ;
        RECT 280.120000 246.260000 281.320000 246.740000 ;
        RECT 280.120000 251.700000 281.320000 252.180000 ;
        RECT 280.120000 257.140000 281.320000 257.620000 ;
        RECT 280.120000 273.460000 281.320000 273.940000 ;
        RECT 280.120000 268.020000 281.320000 268.500000 ;
        RECT 280.120000 262.580000 281.320000 263.060000 ;
        RECT 325.120000 240.820000 326.320000 241.300000 ;
        RECT 325.120000 246.260000 326.320000 246.740000 ;
        RECT 325.120000 251.700000 326.320000 252.180000 ;
        RECT 325.120000 257.140000 326.320000 257.620000 ;
        RECT 325.120000 273.460000 326.320000 273.940000 ;
        RECT 325.120000 268.020000 326.320000 268.500000 ;
        RECT 325.120000 262.580000 326.320000 263.060000 ;
        RECT 370.120000 219.060000 371.320000 219.540000 ;
        RECT 370.120000 213.620000 371.320000 214.100000 ;
        RECT 370.120000 208.180000 371.320000 208.660000 ;
        RECT 370.120000 235.380000 371.320000 235.860000 ;
        RECT 370.120000 224.500000 371.320000 224.980000 ;
        RECT 370.120000 229.940000 371.320000 230.420000 ;
        RECT 370.120000 257.140000 371.320000 257.620000 ;
        RECT 370.120000 251.700000 371.320000 252.180000 ;
        RECT 370.120000 246.260000 371.320000 246.740000 ;
        RECT 370.120000 240.820000 371.320000 241.300000 ;
        RECT 370.120000 273.460000 371.320000 273.940000 ;
        RECT 370.120000 268.020000 371.320000 268.500000 ;
        RECT 370.120000 262.580000 371.320000 263.060000 ;
        RECT 415.120000 137.460000 416.320000 137.940000 ;
        RECT 415.120000 142.900000 416.320000 143.380000 ;
        RECT 415.120000 148.340000 416.320000 148.820000 ;
        RECT 415.120000 153.780000 416.320000 154.260000 ;
        RECT 415.120000 170.100000 416.320000 170.580000 ;
        RECT 415.120000 164.660000 416.320000 165.140000 ;
        RECT 415.120000 159.220000 416.320000 159.700000 ;
        RECT 460.120000 137.460000 461.320000 137.940000 ;
        RECT 460.120000 142.900000 461.320000 143.380000 ;
        RECT 460.120000 148.340000 461.320000 148.820000 ;
        RECT 460.120000 153.780000 461.320000 154.260000 ;
        RECT 460.120000 170.100000 461.320000 170.580000 ;
        RECT 460.120000 164.660000 461.320000 165.140000 ;
        RECT 460.120000 159.220000 461.320000 159.700000 ;
        RECT 415.120000 175.540000 416.320000 176.020000 ;
        RECT 415.120000 180.980000 416.320000 181.460000 ;
        RECT 415.120000 186.420000 416.320000 186.900000 ;
        RECT 415.120000 202.740000 416.320000 203.220000 ;
        RECT 415.120000 197.300000 416.320000 197.780000 ;
        RECT 415.120000 191.860000 416.320000 192.340000 ;
        RECT 460.120000 175.540000 461.320000 176.020000 ;
        RECT 460.120000 180.980000 461.320000 181.460000 ;
        RECT 460.120000 186.420000 461.320000 186.900000 ;
        RECT 460.120000 202.740000 461.320000 203.220000 ;
        RECT 460.120000 197.300000 461.320000 197.780000 ;
        RECT 460.120000 191.860000 461.320000 192.340000 ;
        RECT 505.120000 153.780000 506.320000 154.260000 ;
        RECT 505.120000 148.340000 506.320000 148.820000 ;
        RECT 505.120000 142.900000 506.320000 143.380000 ;
        RECT 505.120000 137.460000 506.320000 137.940000 ;
        RECT 505.120000 170.100000 506.320000 170.580000 ;
        RECT 505.120000 164.660000 506.320000 165.140000 ;
        RECT 505.120000 159.220000 506.320000 159.700000 ;
        RECT 545.600000 153.780000 546.800000 154.260000 ;
        RECT 545.600000 148.340000 546.800000 148.820000 ;
        RECT 545.600000 137.460000 546.800000 137.940000 ;
        RECT 545.600000 142.900000 546.800000 143.380000 ;
        RECT 545.600000 170.100000 546.800000 170.580000 ;
        RECT 545.600000 164.660000 546.800000 165.140000 ;
        RECT 545.600000 159.220000 546.800000 159.700000 ;
        RECT 505.120000 186.420000 506.320000 186.900000 ;
        RECT 505.120000 180.980000 506.320000 181.460000 ;
        RECT 505.120000 175.540000 506.320000 176.020000 ;
        RECT 505.120000 202.740000 506.320000 203.220000 ;
        RECT 505.120000 197.300000 506.320000 197.780000 ;
        RECT 505.120000 191.860000 506.320000 192.340000 ;
        RECT 545.600000 186.420000 546.800000 186.900000 ;
        RECT 545.600000 180.980000 546.800000 181.460000 ;
        RECT 545.600000 175.540000 546.800000 176.020000 ;
        RECT 545.600000 202.740000 546.800000 203.220000 ;
        RECT 545.600000 197.300000 546.800000 197.780000 ;
        RECT 545.600000 191.860000 546.800000 192.340000 ;
        RECT 415.120000 208.180000 416.320000 208.660000 ;
        RECT 415.120000 213.620000 416.320000 214.100000 ;
        RECT 415.120000 219.060000 416.320000 219.540000 ;
        RECT 415.120000 235.380000 416.320000 235.860000 ;
        RECT 415.120000 229.940000 416.320000 230.420000 ;
        RECT 415.120000 224.500000 416.320000 224.980000 ;
        RECT 460.120000 208.180000 461.320000 208.660000 ;
        RECT 460.120000 213.620000 461.320000 214.100000 ;
        RECT 460.120000 219.060000 461.320000 219.540000 ;
        RECT 460.120000 235.380000 461.320000 235.860000 ;
        RECT 460.120000 229.940000 461.320000 230.420000 ;
        RECT 460.120000 224.500000 461.320000 224.980000 ;
        RECT 415.120000 240.820000 416.320000 241.300000 ;
        RECT 415.120000 246.260000 416.320000 246.740000 ;
        RECT 415.120000 251.700000 416.320000 252.180000 ;
        RECT 415.120000 257.140000 416.320000 257.620000 ;
        RECT 415.120000 273.460000 416.320000 273.940000 ;
        RECT 415.120000 268.020000 416.320000 268.500000 ;
        RECT 415.120000 262.580000 416.320000 263.060000 ;
        RECT 460.120000 240.820000 461.320000 241.300000 ;
        RECT 460.120000 246.260000 461.320000 246.740000 ;
        RECT 460.120000 251.700000 461.320000 252.180000 ;
        RECT 460.120000 257.140000 461.320000 257.620000 ;
        RECT 460.120000 273.460000 461.320000 273.940000 ;
        RECT 460.120000 268.020000 461.320000 268.500000 ;
        RECT 460.120000 262.580000 461.320000 263.060000 ;
        RECT 505.120000 219.060000 506.320000 219.540000 ;
        RECT 505.120000 213.620000 506.320000 214.100000 ;
        RECT 505.120000 208.180000 506.320000 208.660000 ;
        RECT 505.120000 235.380000 506.320000 235.860000 ;
        RECT 505.120000 224.500000 506.320000 224.980000 ;
        RECT 505.120000 229.940000 506.320000 230.420000 ;
        RECT 545.600000 219.060000 546.800000 219.540000 ;
        RECT 545.600000 208.180000 546.800000 208.660000 ;
        RECT 545.600000 213.620000 546.800000 214.100000 ;
        RECT 545.600000 235.380000 546.800000 235.860000 ;
        RECT 545.600000 229.940000 546.800000 230.420000 ;
        RECT 545.600000 224.500000 546.800000 224.980000 ;
        RECT 505.120000 257.140000 506.320000 257.620000 ;
        RECT 505.120000 251.700000 506.320000 252.180000 ;
        RECT 505.120000 246.260000 506.320000 246.740000 ;
        RECT 505.120000 240.820000 506.320000 241.300000 ;
        RECT 505.120000 273.460000 506.320000 273.940000 ;
        RECT 505.120000 268.020000 506.320000 268.500000 ;
        RECT 505.120000 262.580000 506.320000 263.060000 ;
        RECT 545.600000 257.140000 546.800000 257.620000 ;
        RECT 545.600000 251.700000 546.800000 252.180000 ;
        RECT 545.600000 240.820000 546.800000 241.300000 ;
        RECT 545.600000 246.260000 546.800000 246.740000 ;
        RECT 545.600000 273.460000 546.800000 273.940000 ;
        RECT 545.600000 268.020000 546.800000 268.500000 ;
        RECT 545.600000 262.580000 546.800000 263.060000 ;
        RECT 3.360000 278.900000 4.560000 279.380000 ;
        RECT 9.955000 278.900000 11.320000 279.380000 ;
        RECT 3.360000 289.780000 4.560000 290.260000 ;
        RECT 9.955000 289.780000 11.320000 290.260000 ;
        RECT 3.360000 284.340000 4.560000 284.820000 ;
        RECT 9.955000 284.340000 11.320000 284.820000 ;
        RECT 3.360000 300.660000 4.560000 301.140000 ;
        RECT 9.955000 300.660000 11.320000 301.140000 ;
        RECT 3.360000 295.220000 4.560000 295.700000 ;
        RECT 9.955000 295.220000 11.320000 295.700000 ;
        RECT 3.360000 306.100000 4.560000 306.580000 ;
        RECT 9.955000 306.100000 11.320000 306.580000 ;
        RECT 55.120000 278.900000 56.320000 279.380000 ;
        RECT 55.120000 284.340000 56.320000 284.820000 ;
        RECT 55.120000 289.780000 56.320000 290.260000 ;
        RECT 55.120000 306.100000 56.320000 306.580000 ;
        RECT 55.120000 300.660000 56.320000 301.140000 ;
        RECT 55.120000 295.220000 56.320000 295.700000 ;
        RECT 3.360000 316.980000 4.560000 317.460000 ;
        RECT 9.955000 316.980000 11.320000 317.460000 ;
        RECT 3.360000 311.540000 4.560000 312.020000 ;
        RECT 9.955000 311.540000 11.320000 312.020000 ;
        RECT 3.360000 322.420000 4.560000 322.900000 ;
        RECT 9.955000 322.420000 11.320000 322.900000 ;
        RECT 3.360000 333.300000 4.560000 333.780000 ;
        RECT 9.955000 333.300000 11.320000 333.780000 ;
        RECT 3.360000 327.860000 4.560000 328.340000 ;
        RECT 9.955000 327.860000 11.320000 328.340000 ;
        RECT 3.360000 338.740000 4.560000 339.220000 ;
        RECT 9.955000 338.740000 11.320000 339.220000 ;
        RECT 55.120000 311.540000 56.320000 312.020000 ;
        RECT 55.120000 316.980000 56.320000 317.460000 ;
        RECT 55.120000 322.420000 56.320000 322.900000 ;
        RECT 55.120000 338.740000 56.320000 339.220000 ;
        RECT 55.120000 333.300000 56.320000 333.780000 ;
        RECT 55.120000 327.860000 56.320000 328.340000 ;
        RECT 100.120000 306.100000 101.320000 306.580000 ;
        RECT 100.120000 300.660000 101.320000 301.140000 ;
        RECT 100.120000 278.900000 101.320000 279.380000 ;
        RECT 100.120000 284.340000 101.320000 284.820000 ;
        RECT 100.120000 289.780000 101.320000 290.260000 ;
        RECT 100.120000 295.220000 101.320000 295.700000 ;
        RECT 100.120000 338.740000 101.320000 339.220000 ;
        RECT 100.120000 333.300000 101.320000 333.780000 ;
        RECT 100.120000 311.540000 101.320000 312.020000 ;
        RECT 100.120000 316.980000 101.320000 317.460000 ;
        RECT 100.120000 322.420000 101.320000 322.900000 ;
        RECT 100.120000 327.860000 101.320000 328.340000 ;
        RECT 3.360000 360.500000 4.560000 360.980000 ;
        RECT 9.955000 360.500000 11.320000 360.980000 ;
        RECT 3.360000 349.620000 4.560000 350.100000 ;
        RECT 9.955000 349.620000 11.320000 350.100000 ;
        RECT 3.360000 344.180000 4.560000 344.660000 ;
        RECT 9.955000 344.180000 11.320000 344.660000 ;
        RECT 3.360000 355.060000 4.560000 355.540000 ;
        RECT 9.955000 355.060000 11.320000 355.540000 ;
        RECT 3.360000 365.940000 4.560000 366.420000 ;
        RECT 9.955000 365.940000 11.320000 366.420000 ;
        RECT 3.360000 376.820000 4.560000 377.300000 ;
        RECT 9.955000 376.820000 11.320000 377.300000 ;
        RECT 3.360000 371.380000 4.560000 371.860000 ;
        RECT 9.955000 371.380000 11.320000 371.860000 ;
        RECT 55.120000 360.500000 56.320000 360.980000 ;
        RECT 55.120000 344.180000 56.320000 344.660000 ;
        RECT 55.120000 349.620000 56.320000 350.100000 ;
        RECT 55.120000 355.060000 56.320000 355.540000 ;
        RECT 55.120000 376.820000 56.320000 377.300000 ;
        RECT 55.120000 371.380000 56.320000 371.860000 ;
        RECT 55.120000 365.940000 56.320000 366.420000 ;
        RECT 3.360000 382.260000 4.560000 382.740000 ;
        RECT 9.955000 382.260000 11.320000 382.740000 ;
        RECT 3.360000 393.140000 4.560000 393.620000 ;
        RECT 9.955000 393.140000 11.320000 393.620000 ;
        RECT 3.360000 387.700000 4.560000 388.180000 ;
        RECT 9.955000 387.700000 11.320000 388.180000 ;
        RECT 3.360000 398.580000 4.560000 399.060000 ;
        RECT 9.955000 398.580000 11.320000 399.060000 ;
        RECT 3.360000 409.460000 4.560000 409.940000 ;
        RECT 9.955000 409.460000 11.320000 409.940000 ;
        RECT 3.360000 404.020000 4.560000 404.500000 ;
        RECT 9.955000 404.020000 11.320000 404.500000 ;
        RECT 55.120000 382.260000 56.320000 382.740000 ;
        RECT 55.120000 387.700000 56.320000 388.180000 ;
        RECT 55.120000 393.140000 56.320000 393.620000 ;
        RECT 55.120000 409.460000 56.320000 409.940000 ;
        RECT 55.120000 404.020000 56.320000 404.500000 ;
        RECT 55.120000 398.580000 56.320000 399.060000 ;
        RECT 100.120000 376.820000 101.320000 377.300000 ;
        RECT 100.120000 371.380000 101.320000 371.860000 ;
        RECT 100.120000 365.940000 101.320000 366.420000 ;
        RECT 100.120000 344.180000 101.320000 344.660000 ;
        RECT 100.120000 349.620000 101.320000 350.100000 ;
        RECT 100.120000 355.060000 101.320000 355.540000 ;
        RECT 100.120000 360.500000 101.320000 360.980000 ;
        RECT 100.120000 409.460000 101.320000 409.940000 ;
        RECT 100.120000 404.020000 101.320000 404.500000 ;
        RECT 100.120000 382.260000 101.320000 382.740000 ;
        RECT 100.120000 387.700000 101.320000 388.180000 ;
        RECT 100.120000 393.140000 101.320000 393.620000 ;
        RECT 100.120000 398.580000 101.320000 399.060000 ;
        RECT 145.120000 278.900000 146.320000 279.380000 ;
        RECT 145.120000 284.340000 146.320000 284.820000 ;
        RECT 145.120000 289.780000 146.320000 290.260000 ;
        RECT 145.120000 306.100000 146.320000 306.580000 ;
        RECT 145.120000 300.660000 146.320000 301.140000 ;
        RECT 145.120000 295.220000 146.320000 295.700000 ;
        RECT 190.120000 278.900000 191.320000 279.380000 ;
        RECT 190.120000 284.340000 191.320000 284.820000 ;
        RECT 190.120000 289.780000 191.320000 290.260000 ;
        RECT 190.120000 306.100000 191.320000 306.580000 ;
        RECT 190.120000 300.660000 191.320000 301.140000 ;
        RECT 190.120000 295.220000 191.320000 295.700000 ;
        RECT 145.120000 311.540000 146.320000 312.020000 ;
        RECT 145.120000 316.980000 146.320000 317.460000 ;
        RECT 145.120000 322.420000 146.320000 322.900000 ;
        RECT 145.120000 338.740000 146.320000 339.220000 ;
        RECT 145.120000 333.300000 146.320000 333.780000 ;
        RECT 145.120000 327.860000 146.320000 328.340000 ;
        RECT 190.120000 311.540000 191.320000 312.020000 ;
        RECT 190.120000 316.980000 191.320000 317.460000 ;
        RECT 190.120000 322.420000 191.320000 322.900000 ;
        RECT 190.120000 338.740000 191.320000 339.220000 ;
        RECT 190.120000 333.300000 191.320000 333.780000 ;
        RECT 190.120000 327.860000 191.320000 328.340000 ;
        RECT 235.120000 289.780000 236.320000 290.260000 ;
        RECT 235.120000 284.340000 236.320000 284.820000 ;
        RECT 235.120000 278.900000 236.320000 279.380000 ;
        RECT 235.120000 306.100000 236.320000 306.580000 ;
        RECT 235.120000 295.220000 236.320000 295.700000 ;
        RECT 235.120000 300.660000 236.320000 301.140000 ;
        RECT 235.120000 322.420000 236.320000 322.900000 ;
        RECT 235.120000 316.980000 236.320000 317.460000 ;
        RECT 235.120000 311.540000 236.320000 312.020000 ;
        RECT 235.120000 338.740000 236.320000 339.220000 ;
        RECT 235.120000 327.860000 236.320000 328.340000 ;
        RECT 235.120000 333.300000 236.320000 333.780000 ;
        RECT 145.120000 360.500000 146.320000 360.980000 ;
        RECT 145.120000 344.180000 146.320000 344.660000 ;
        RECT 145.120000 349.620000 146.320000 350.100000 ;
        RECT 145.120000 355.060000 146.320000 355.540000 ;
        RECT 145.120000 376.820000 146.320000 377.300000 ;
        RECT 145.120000 371.380000 146.320000 371.860000 ;
        RECT 145.120000 365.940000 146.320000 366.420000 ;
        RECT 190.120000 360.500000 191.320000 360.980000 ;
        RECT 190.120000 344.180000 191.320000 344.660000 ;
        RECT 190.120000 349.620000 191.320000 350.100000 ;
        RECT 190.120000 355.060000 191.320000 355.540000 ;
        RECT 190.120000 376.820000 191.320000 377.300000 ;
        RECT 190.120000 371.380000 191.320000 371.860000 ;
        RECT 190.120000 365.940000 191.320000 366.420000 ;
        RECT 145.120000 382.260000 146.320000 382.740000 ;
        RECT 145.120000 387.700000 146.320000 388.180000 ;
        RECT 145.120000 393.140000 146.320000 393.620000 ;
        RECT 145.120000 409.460000 146.320000 409.940000 ;
        RECT 145.120000 404.020000 146.320000 404.500000 ;
        RECT 145.120000 398.580000 146.320000 399.060000 ;
        RECT 190.120000 382.260000 191.320000 382.740000 ;
        RECT 190.120000 387.700000 191.320000 388.180000 ;
        RECT 190.120000 393.140000 191.320000 393.620000 ;
        RECT 190.120000 409.460000 191.320000 409.940000 ;
        RECT 190.120000 404.020000 191.320000 404.500000 ;
        RECT 190.120000 398.580000 191.320000 399.060000 ;
        RECT 235.120000 360.500000 236.320000 360.980000 ;
        RECT 235.120000 355.060000 236.320000 355.540000 ;
        RECT 235.120000 349.620000 236.320000 350.100000 ;
        RECT 235.120000 344.180000 236.320000 344.660000 ;
        RECT 235.120000 376.820000 236.320000 377.300000 ;
        RECT 235.120000 371.380000 236.320000 371.860000 ;
        RECT 235.120000 365.940000 236.320000 366.420000 ;
        RECT 235.120000 393.140000 236.320000 393.620000 ;
        RECT 235.120000 387.700000 236.320000 388.180000 ;
        RECT 235.120000 382.260000 236.320000 382.740000 ;
        RECT 235.120000 409.460000 236.320000 409.940000 ;
        RECT 235.120000 398.580000 236.320000 399.060000 ;
        RECT 235.120000 404.020000 236.320000 404.500000 ;
        RECT 3.360000 420.340000 4.560000 420.820000 ;
        RECT 9.955000 420.340000 11.320000 420.820000 ;
        RECT 3.360000 414.900000 4.560000 415.380000 ;
        RECT 9.955000 414.900000 11.320000 415.380000 ;
        RECT 3.360000 425.780000 4.560000 426.260000 ;
        RECT 9.955000 425.780000 11.320000 426.260000 ;
        RECT 3.360000 436.660000 4.560000 437.140000 ;
        RECT 9.955000 436.660000 11.320000 437.140000 ;
        RECT 3.360000 431.220000 4.560000 431.700000 ;
        RECT 9.955000 431.220000 11.320000 431.700000 ;
        RECT 3.360000 442.100000 4.560000 442.580000 ;
        RECT 9.955000 442.100000 11.320000 442.580000 ;
        RECT 55.120000 414.900000 56.320000 415.380000 ;
        RECT 55.120000 420.340000 56.320000 420.820000 ;
        RECT 55.120000 425.780000 56.320000 426.260000 ;
        RECT 55.120000 442.100000 56.320000 442.580000 ;
        RECT 55.120000 436.660000 56.320000 437.140000 ;
        RECT 55.120000 431.220000 56.320000 431.700000 ;
        RECT 3.360000 463.860000 4.560000 464.340000 ;
        RECT 9.955000 463.860000 11.320000 464.340000 ;
        RECT 3.360000 452.980000 4.560000 453.460000 ;
        RECT 9.955000 452.980000 11.320000 453.460000 ;
        RECT 3.360000 447.540000 4.560000 448.020000 ;
        RECT 9.955000 447.540000 11.320000 448.020000 ;
        RECT 3.360000 458.420000 4.560000 458.900000 ;
        RECT 9.955000 458.420000 11.320000 458.900000 ;
        RECT 3.360000 469.300000 4.560000 469.780000 ;
        RECT 9.955000 469.300000 11.320000 469.780000 ;
        RECT 3.360000 480.180000 4.560000 480.660000 ;
        RECT 9.955000 480.180000 11.320000 480.660000 ;
        RECT 3.360000 474.740000 4.560000 475.220000 ;
        RECT 9.955000 474.740000 11.320000 475.220000 ;
        RECT 55.120000 463.860000 56.320000 464.340000 ;
        RECT 55.120000 447.540000 56.320000 448.020000 ;
        RECT 55.120000 452.980000 56.320000 453.460000 ;
        RECT 55.120000 458.420000 56.320000 458.900000 ;
        RECT 55.120000 480.180000 56.320000 480.660000 ;
        RECT 55.120000 474.740000 56.320000 475.220000 ;
        RECT 55.120000 469.300000 56.320000 469.780000 ;
        RECT 100.120000 442.100000 101.320000 442.580000 ;
        RECT 100.120000 436.660000 101.320000 437.140000 ;
        RECT 100.120000 414.900000 101.320000 415.380000 ;
        RECT 100.120000 420.340000 101.320000 420.820000 ;
        RECT 100.120000 425.780000 101.320000 426.260000 ;
        RECT 100.120000 431.220000 101.320000 431.700000 ;
        RECT 100.120000 480.180000 101.320000 480.660000 ;
        RECT 100.120000 474.740000 101.320000 475.220000 ;
        RECT 100.120000 469.300000 101.320000 469.780000 ;
        RECT 100.120000 447.540000 101.320000 448.020000 ;
        RECT 100.120000 452.980000 101.320000 453.460000 ;
        RECT 100.120000 458.420000 101.320000 458.900000 ;
        RECT 100.120000 463.860000 101.320000 464.340000 ;
        RECT 3.360000 485.620000 4.560000 486.100000 ;
        RECT 9.955000 485.620000 11.320000 486.100000 ;
        RECT 3.360000 496.500000 4.560000 496.980000 ;
        RECT 9.955000 496.500000 11.320000 496.980000 ;
        RECT 3.360000 491.060000 4.560000 491.540000 ;
        RECT 9.955000 491.060000 11.320000 491.540000 ;
        RECT 3.360000 501.940000 4.560000 502.420000 ;
        RECT 9.955000 501.940000 11.320000 502.420000 ;
        RECT 3.360000 512.820000 4.560000 513.300000 ;
        RECT 9.955000 512.820000 11.320000 513.300000 ;
        RECT 3.360000 507.380000 4.560000 507.860000 ;
        RECT 9.955000 507.380000 11.320000 507.860000 ;
        RECT 55.120000 485.620000 56.320000 486.100000 ;
        RECT 55.120000 491.060000 56.320000 491.540000 ;
        RECT 55.120000 496.500000 56.320000 496.980000 ;
        RECT 55.120000 512.820000 56.320000 513.300000 ;
        RECT 55.120000 507.380000 56.320000 507.860000 ;
        RECT 55.120000 501.940000 56.320000 502.420000 ;
        RECT 3.360000 523.700000 4.560000 524.180000 ;
        RECT 9.955000 523.700000 11.320000 524.180000 ;
        RECT 3.360000 518.260000 4.560000 518.740000 ;
        RECT 9.955000 518.260000 11.320000 518.740000 ;
        RECT 3.360000 529.140000 4.560000 529.620000 ;
        RECT 9.955000 529.140000 11.320000 529.620000 ;
        RECT 3.360000 534.580000 4.560000 535.060000 ;
        RECT 9.955000 534.580000 11.320000 535.060000 ;
        RECT 55.120000 534.580000 56.320000 535.060000 ;
        RECT 55.120000 529.140000 56.320000 529.620000 ;
        RECT 55.120000 523.700000 56.320000 524.180000 ;
        RECT 55.120000 518.260000 56.320000 518.740000 ;
        RECT 100.120000 512.820000 101.320000 513.300000 ;
        RECT 100.120000 507.380000 101.320000 507.860000 ;
        RECT 100.120000 485.620000 101.320000 486.100000 ;
        RECT 100.120000 491.060000 101.320000 491.540000 ;
        RECT 100.120000 496.500000 101.320000 496.980000 ;
        RECT 100.120000 501.940000 101.320000 502.420000 ;
        RECT 100.120000 534.580000 101.320000 535.060000 ;
        RECT 100.120000 529.140000 101.320000 529.620000 ;
        RECT 100.120000 523.700000 101.320000 524.180000 ;
        RECT 100.120000 518.260000 101.320000 518.740000 ;
        RECT 145.120000 414.900000 146.320000 415.380000 ;
        RECT 145.120000 420.340000 146.320000 420.820000 ;
        RECT 145.120000 425.780000 146.320000 426.260000 ;
        RECT 145.120000 442.100000 146.320000 442.580000 ;
        RECT 145.120000 436.660000 146.320000 437.140000 ;
        RECT 145.120000 431.220000 146.320000 431.700000 ;
        RECT 190.120000 414.900000 191.320000 415.380000 ;
        RECT 190.120000 420.340000 191.320000 420.820000 ;
        RECT 190.120000 425.780000 191.320000 426.260000 ;
        RECT 190.120000 442.100000 191.320000 442.580000 ;
        RECT 190.120000 436.660000 191.320000 437.140000 ;
        RECT 190.120000 431.220000 191.320000 431.700000 ;
        RECT 145.120000 463.860000 146.320000 464.340000 ;
        RECT 145.120000 447.540000 146.320000 448.020000 ;
        RECT 145.120000 452.980000 146.320000 453.460000 ;
        RECT 145.120000 458.420000 146.320000 458.900000 ;
        RECT 145.120000 480.180000 146.320000 480.660000 ;
        RECT 145.120000 474.740000 146.320000 475.220000 ;
        RECT 145.120000 469.300000 146.320000 469.780000 ;
        RECT 190.120000 463.860000 191.320000 464.340000 ;
        RECT 190.120000 447.540000 191.320000 448.020000 ;
        RECT 190.120000 452.980000 191.320000 453.460000 ;
        RECT 190.120000 458.420000 191.320000 458.900000 ;
        RECT 190.120000 480.180000 191.320000 480.660000 ;
        RECT 190.120000 474.740000 191.320000 475.220000 ;
        RECT 190.120000 469.300000 191.320000 469.780000 ;
        RECT 235.120000 425.780000 236.320000 426.260000 ;
        RECT 235.120000 420.340000 236.320000 420.820000 ;
        RECT 235.120000 414.900000 236.320000 415.380000 ;
        RECT 235.120000 442.100000 236.320000 442.580000 ;
        RECT 235.120000 431.220000 236.320000 431.700000 ;
        RECT 235.120000 436.660000 236.320000 437.140000 ;
        RECT 235.120000 463.860000 236.320000 464.340000 ;
        RECT 235.120000 458.420000 236.320000 458.900000 ;
        RECT 235.120000 452.980000 236.320000 453.460000 ;
        RECT 235.120000 447.540000 236.320000 448.020000 ;
        RECT 235.120000 480.180000 236.320000 480.660000 ;
        RECT 235.120000 474.740000 236.320000 475.220000 ;
        RECT 235.120000 469.300000 236.320000 469.780000 ;
        RECT 145.120000 485.620000 146.320000 486.100000 ;
        RECT 145.120000 491.060000 146.320000 491.540000 ;
        RECT 145.120000 496.500000 146.320000 496.980000 ;
        RECT 145.120000 512.820000 146.320000 513.300000 ;
        RECT 145.120000 507.380000 146.320000 507.860000 ;
        RECT 145.120000 501.940000 146.320000 502.420000 ;
        RECT 190.120000 485.620000 191.320000 486.100000 ;
        RECT 190.120000 491.060000 191.320000 491.540000 ;
        RECT 190.120000 496.500000 191.320000 496.980000 ;
        RECT 190.120000 512.820000 191.320000 513.300000 ;
        RECT 190.120000 507.380000 191.320000 507.860000 ;
        RECT 190.120000 501.940000 191.320000 502.420000 ;
        RECT 145.120000 534.580000 146.320000 535.060000 ;
        RECT 145.120000 529.140000 146.320000 529.620000 ;
        RECT 145.120000 523.700000 146.320000 524.180000 ;
        RECT 145.120000 518.260000 146.320000 518.740000 ;
        RECT 190.120000 534.580000 191.320000 535.060000 ;
        RECT 190.120000 529.140000 191.320000 529.620000 ;
        RECT 190.120000 523.700000 191.320000 524.180000 ;
        RECT 190.120000 518.260000 191.320000 518.740000 ;
        RECT 235.120000 496.500000 236.320000 496.980000 ;
        RECT 235.120000 491.060000 236.320000 491.540000 ;
        RECT 235.120000 485.620000 236.320000 486.100000 ;
        RECT 235.120000 512.820000 236.320000 513.300000 ;
        RECT 235.120000 501.940000 236.320000 502.420000 ;
        RECT 235.120000 507.380000 236.320000 507.860000 ;
        RECT 235.120000 534.580000 236.320000 535.060000 ;
        RECT 235.120000 529.140000 236.320000 529.620000 ;
        RECT 235.120000 523.700000 236.320000 524.180000 ;
        RECT 235.120000 518.260000 236.320000 518.740000 ;
        RECT 280.120000 278.900000 281.320000 279.380000 ;
        RECT 280.120000 284.340000 281.320000 284.820000 ;
        RECT 280.120000 289.780000 281.320000 290.260000 ;
        RECT 280.120000 306.100000 281.320000 306.580000 ;
        RECT 280.120000 300.660000 281.320000 301.140000 ;
        RECT 280.120000 295.220000 281.320000 295.700000 ;
        RECT 325.120000 278.900000 326.320000 279.380000 ;
        RECT 325.120000 284.340000 326.320000 284.820000 ;
        RECT 325.120000 289.780000 326.320000 290.260000 ;
        RECT 325.120000 306.100000 326.320000 306.580000 ;
        RECT 325.120000 300.660000 326.320000 301.140000 ;
        RECT 325.120000 295.220000 326.320000 295.700000 ;
        RECT 280.120000 311.540000 281.320000 312.020000 ;
        RECT 280.120000 316.980000 281.320000 317.460000 ;
        RECT 280.120000 322.420000 281.320000 322.900000 ;
        RECT 280.120000 338.740000 281.320000 339.220000 ;
        RECT 280.120000 333.300000 281.320000 333.780000 ;
        RECT 280.120000 327.860000 281.320000 328.340000 ;
        RECT 325.120000 311.540000 326.320000 312.020000 ;
        RECT 325.120000 316.980000 326.320000 317.460000 ;
        RECT 325.120000 322.420000 326.320000 322.900000 ;
        RECT 325.120000 338.740000 326.320000 339.220000 ;
        RECT 325.120000 333.300000 326.320000 333.780000 ;
        RECT 325.120000 327.860000 326.320000 328.340000 ;
        RECT 370.120000 289.780000 371.320000 290.260000 ;
        RECT 370.120000 284.340000 371.320000 284.820000 ;
        RECT 370.120000 278.900000 371.320000 279.380000 ;
        RECT 370.120000 306.100000 371.320000 306.580000 ;
        RECT 370.120000 295.220000 371.320000 295.700000 ;
        RECT 370.120000 300.660000 371.320000 301.140000 ;
        RECT 370.120000 322.420000 371.320000 322.900000 ;
        RECT 370.120000 316.980000 371.320000 317.460000 ;
        RECT 370.120000 311.540000 371.320000 312.020000 ;
        RECT 370.120000 338.740000 371.320000 339.220000 ;
        RECT 370.120000 327.860000 371.320000 328.340000 ;
        RECT 370.120000 333.300000 371.320000 333.780000 ;
        RECT 280.120000 360.500000 281.320000 360.980000 ;
        RECT 280.120000 344.180000 281.320000 344.660000 ;
        RECT 280.120000 349.620000 281.320000 350.100000 ;
        RECT 280.120000 355.060000 281.320000 355.540000 ;
        RECT 280.120000 376.820000 281.320000 377.300000 ;
        RECT 280.120000 371.380000 281.320000 371.860000 ;
        RECT 280.120000 365.940000 281.320000 366.420000 ;
        RECT 325.120000 360.500000 326.320000 360.980000 ;
        RECT 325.120000 344.180000 326.320000 344.660000 ;
        RECT 325.120000 349.620000 326.320000 350.100000 ;
        RECT 325.120000 355.060000 326.320000 355.540000 ;
        RECT 325.120000 376.820000 326.320000 377.300000 ;
        RECT 325.120000 371.380000 326.320000 371.860000 ;
        RECT 325.120000 365.940000 326.320000 366.420000 ;
        RECT 280.120000 382.260000 281.320000 382.740000 ;
        RECT 280.120000 387.700000 281.320000 388.180000 ;
        RECT 280.120000 393.140000 281.320000 393.620000 ;
        RECT 280.120000 409.460000 281.320000 409.940000 ;
        RECT 280.120000 404.020000 281.320000 404.500000 ;
        RECT 280.120000 398.580000 281.320000 399.060000 ;
        RECT 325.120000 382.260000 326.320000 382.740000 ;
        RECT 325.120000 387.700000 326.320000 388.180000 ;
        RECT 325.120000 393.140000 326.320000 393.620000 ;
        RECT 325.120000 409.460000 326.320000 409.940000 ;
        RECT 325.120000 404.020000 326.320000 404.500000 ;
        RECT 325.120000 398.580000 326.320000 399.060000 ;
        RECT 370.120000 360.500000 371.320000 360.980000 ;
        RECT 370.120000 355.060000 371.320000 355.540000 ;
        RECT 370.120000 349.620000 371.320000 350.100000 ;
        RECT 370.120000 344.180000 371.320000 344.660000 ;
        RECT 370.120000 376.820000 371.320000 377.300000 ;
        RECT 370.120000 371.380000 371.320000 371.860000 ;
        RECT 370.120000 365.940000 371.320000 366.420000 ;
        RECT 370.120000 393.140000 371.320000 393.620000 ;
        RECT 370.120000 387.700000 371.320000 388.180000 ;
        RECT 370.120000 382.260000 371.320000 382.740000 ;
        RECT 370.120000 409.460000 371.320000 409.940000 ;
        RECT 370.120000 398.580000 371.320000 399.060000 ;
        RECT 370.120000 404.020000 371.320000 404.500000 ;
        RECT 415.120000 278.900000 416.320000 279.380000 ;
        RECT 415.120000 284.340000 416.320000 284.820000 ;
        RECT 415.120000 289.780000 416.320000 290.260000 ;
        RECT 415.120000 306.100000 416.320000 306.580000 ;
        RECT 415.120000 300.660000 416.320000 301.140000 ;
        RECT 415.120000 295.220000 416.320000 295.700000 ;
        RECT 460.120000 278.900000 461.320000 279.380000 ;
        RECT 460.120000 284.340000 461.320000 284.820000 ;
        RECT 460.120000 289.780000 461.320000 290.260000 ;
        RECT 460.120000 306.100000 461.320000 306.580000 ;
        RECT 460.120000 300.660000 461.320000 301.140000 ;
        RECT 460.120000 295.220000 461.320000 295.700000 ;
        RECT 415.120000 311.540000 416.320000 312.020000 ;
        RECT 415.120000 316.980000 416.320000 317.460000 ;
        RECT 415.120000 322.420000 416.320000 322.900000 ;
        RECT 415.120000 338.740000 416.320000 339.220000 ;
        RECT 415.120000 333.300000 416.320000 333.780000 ;
        RECT 415.120000 327.860000 416.320000 328.340000 ;
        RECT 460.120000 311.540000 461.320000 312.020000 ;
        RECT 460.120000 316.980000 461.320000 317.460000 ;
        RECT 460.120000 322.420000 461.320000 322.900000 ;
        RECT 460.120000 338.740000 461.320000 339.220000 ;
        RECT 460.120000 333.300000 461.320000 333.780000 ;
        RECT 460.120000 327.860000 461.320000 328.340000 ;
        RECT 505.120000 289.780000 506.320000 290.260000 ;
        RECT 505.120000 284.340000 506.320000 284.820000 ;
        RECT 505.120000 278.900000 506.320000 279.380000 ;
        RECT 505.120000 306.100000 506.320000 306.580000 ;
        RECT 505.120000 295.220000 506.320000 295.700000 ;
        RECT 505.120000 300.660000 506.320000 301.140000 ;
        RECT 545.600000 289.780000 546.800000 290.260000 ;
        RECT 545.600000 278.900000 546.800000 279.380000 ;
        RECT 545.600000 284.340000 546.800000 284.820000 ;
        RECT 545.600000 306.100000 546.800000 306.580000 ;
        RECT 545.600000 300.660000 546.800000 301.140000 ;
        RECT 545.600000 295.220000 546.800000 295.700000 ;
        RECT 505.120000 322.420000 506.320000 322.900000 ;
        RECT 505.120000 316.980000 506.320000 317.460000 ;
        RECT 505.120000 311.540000 506.320000 312.020000 ;
        RECT 505.120000 338.740000 506.320000 339.220000 ;
        RECT 505.120000 327.860000 506.320000 328.340000 ;
        RECT 505.120000 333.300000 506.320000 333.780000 ;
        RECT 545.600000 322.420000 546.800000 322.900000 ;
        RECT 545.600000 311.540000 546.800000 312.020000 ;
        RECT 545.600000 316.980000 546.800000 317.460000 ;
        RECT 545.600000 338.740000 546.800000 339.220000 ;
        RECT 545.600000 333.300000 546.800000 333.780000 ;
        RECT 545.600000 327.860000 546.800000 328.340000 ;
        RECT 415.120000 360.500000 416.320000 360.980000 ;
        RECT 415.120000 344.180000 416.320000 344.660000 ;
        RECT 415.120000 349.620000 416.320000 350.100000 ;
        RECT 415.120000 355.060000 416.320000 355.540000 ;
        RECT 415.120000 376.820000 416.320000 377.300000 ;
        RECT 415.120000 371.380000 416.320000 371.860000 ;
        RECT 415.120000 365.940000 416.320000 366.420000 ;
        RECT 460.120000 360.500000 461.320000 360.980000 ;
        RECT 460.120000 344.180000 461.320000 344.660000 ;
        RECT 460.120000 349.620000 461.320000 350.100000 ;
        RECT 460.120000 355.060000 461.320000 355.540000 ;
        RECT 460.120000 376.820000 461.320000 377.300000 ;
        RECT 460.120000 371.380000 461.320000 371.860000 ;
        RECT 460.120000 365.940000 461.320000 366.420000 ;
        RECT 415.120000 382.260000 416.320000 382.740000 ;
        RECT 415.120000 387.700000 416.320000 388.180000 ;
        RECT 415.120000 393.140000 416.320000 393.620000 ;
        RECT 415.120000 409.460000 416.320000 409.940000 ;
        RECT 415.120000 404.020000 416.320000 404.500000 ;
        RECT 415.120000 398.580000 416.320000 399.060000 ;
        RECT 460.120000 382.260000 461.320000 382.740000 ;
        RECT 460.120000 387.700000 461.320000 388.180000 ;
        RECT 460.120000 393.140000 461.320000 393.620000 ;
        RECT 460.120000 409.460000 461.320000 409.940000 ;
        RECT 460.120000 404.020000 461.320000 404.500000 ;
        RECT 460.120000 398.580000 461.320000 399.060000 ;
        RECT 505.120000 360.500000 506.320000 360.980000 ;
        RECT 505.120000 355.060000 506.320000 355.540000 ;
        RECT 505.120000 349.620000 506.320000 350.100000 ;
        RECT 505.120000 344.180000 506.320000 344.660000 ;
        RECT 505.120000 376.820000 506.320000 377.300000 ;
        RECT 505.120000 371.380000 506.320000 371.860000 ;
        RECT 505.120000 365.940000 506.320000 366.420000 ;
        RECT 545.600000 360.500000 546.800000 360.980000 ;
        RECT 545.600000 355.060000 546.800000 355.540000 ;
        RECT 545.600000 344.180000 546.800000 344.660000 ;
        RECT 545.600000 349.620000 546.800000 350.100000 ;
        RECT 545.600000 376.820000 546.800000 377.300000 ;
        RECT 545.600000 371.380000 546.800000 371.860000 ;
        RECT 545.600000 365.940000 546.800000 366.420000 ;
        RECT 505.120000 393.140000 506.320000 393.620000 ;
        RECT 505.120000 387.700000 506.320000 388.180000 ;
        RECT 505.120000 382.260000 506.320000 382.740000 ;
        RECT 505.120000 409.460000 506.320000 409.940000 ;
        RECT 505.120000 398.580000 506.320000 399.060000 ;
        RECT 505.120000 404.020000 506.320000 404.500000 ;
        RECT 545.600000 393.140000 546.800000 393.620000 ;
        RECT 545.600000 382.260000 546.800000 382.740000 ;
        RECT 545.600000 387.700000 546.800000 388.180000 ;
        RECT 545.600000 409.460000 546.800000 409.940000 ;
        RECT 545.600000 404.020000 546.800000 404.500000 ;
        RECT 545.600000 398.580000 546.800000 399.060000 ;
        RECT 280.120000 414.900000 281.320000 415.380000 ;
        RECT 280.120000 420.340000 281.320000 420.820000 ;
        RECT 280.120000 425.780000 281.320000 426.260000 ;
        RECT 280.120000 442.100000 281.320000 442.580000 ;
        RECT 280.120000 436.660000 281.320000 437.140000 ;
        RECT 280.120000 431.220000 281.320000 431.700000 ;
        RECT 325.120000 414.900000 326.320000 415.380000 ;
        RECT 325.120000 420.340000 326.320000 420.820000 ;
        RECT 325.120000 425.780000 326.320000 426.260000 ;
        RECT 325.120000 442.100000 326.320000 442.580000 ;
        RECT 325.120000 436.660000 326.320000 437.140000 ;
        RECT 325.120000 431.220000 326.320000 431.700000 ;
        RECT 280.120000 463.860000 281.320000 464.340000 ;
        RECT 280.120000 447.540000 281.320000 448.020000 ;
        RECT 280.120000 452.980000 281.320000 453.460000 ;
        RECT 280.120000 458.420000 281.320000 458.900000 ;
        RECT 280.120000 480.180000 281.320000 480.660000 ;
        RECT 280.120000 474.740000 281.320000 475.220000 ;
        RECT 280.120000 469.300000 281.320000 469.780000 ;
        RECT 325.120000 463.860000 326.320000 464.340000 ;
        RECT 325.120000 447.540000 326.320000 448.020000 ;
        RECT 325.120000 452.980000 326.320000 453.460000 ;
        RECT 325.120000 458.420000 326.320000 458.900000 ;
        RECT 325.120000 480.180000 326.320000 480.660000 ;
        RECT 325.120000 474.740000 326.320000 475.220000 ;
        RECT 325.120000 469.300000 326.320000 469.780000 ;
        RECT 370.120000 425.780000 371.320000 426.260000 ;
        RECT 370.120000 420.340000 371.320000 420.820000 ;
        RECT 370.120000 414.900000 371.320000 415.380000 ;
        RECT 370.120000 442.100000 371.320000 442.580000 ;
        RECT 370.120000 431.220000 371.320000 431.700000 ;
        RECT 370.120000 436.660000 371.320000 437.140000 ;
        RECT 370.120000 463.860000 371.320000 464.340000 ;
        RECT 370.120000 458.420000 371.320000 458.900000 ;
        RECT 370.120000 452.980000 371.320000 453.460000 ;
        RECT 370.120000 447.540000 371.320000 448.020000 ;
        RECT 370.120000 480.180000 371.320000 480.660000 ;
        RECT 370.120000 474.740000 371.320000 475.220000 ;
        RECT 370.120000 469.300000 371.320000 469.780000 ;
        RECT 280.120000 485.620000 281.320000 486.100000 ;
        RECT 280.120000 491.060000 281.320000 491.540000 ;
        RECT 280.120000 496.500000 281.320000 496.980000 ;
        RECT 280.120000 512.820000 281.320000 513.300000 ;
        RECT 280.120000 507.380000 281.320000 507.860000 ;
        RECT 280.120000 501.940000 281.320000 502.420000 ;
        RECT 325.120000 485.620000 326.320000 486.100000 ;
        RECT 325.120000 491.060000 326.320000 491.540000 ;
        RECT 325.120000 496.500000 326.320000 496.980000 ;
        RECT 325.120000 512.820000 326.320000 513.300000 ;
        RECT 325.120000 507.380000 326.320000 507.860000 ;
        RECT 325.120000 501.940000 326.320000 502.420000 ;
        RECT 280.120000 534.580000 281.320000 535.060000 ;
        RECT 280.120000 529.140000 281.320000 529.620000 ;
        RECT 280.120000 523.700000 281.320000 524.180000 ;
        RECT 280.120000 518.260000 281.320000 518.740000 ;
        RECT 325.120000 534.580000 326.320000 535.060000 ;
        RECT 325.120000 529.140000 326.320000 529.620000 ;
        RECT 325.120000 523.700000 326.320000 524.180000 ;
        RECT 325.120000 518.260000 326.320000 518.740000 ;
        RECT 370.120000 496.500000 371.320000 496.980000 ;
        RECT 370.120000 491.060000 371.320000 491.540000 ;
        RECT 370.120000 485.620000 371.320000 486.100000 ;
        RECT 370.120000 512.820000 371.320000 513.300000 ;
        RECT 370.120000 501.940000 371.320000 502.420000 ;
        RECT 370.120000 507.380000 371.320000 507.860000 ;
        RECT 370.120000 534.580000 371.320000 535.060000 ;
        RECT 370.120000 529.140000 371.320000 529.620000 ;
        RECT 370.120000 523.700000 371.320000 524.180000 ;
        RECT 370.120000 518.260000 371.320000 518.740000 ;
        RECT 415.120000 414.900000 416.320000 415.380000 ;
        RECT 415.120000 420.340000 416.320000 420.820000 ;
        RECT 415.120000 425.780000 416.320000 426.260000 ;
        RECT 415.120000 442.100000 416.320000 442.580000 ;
        RECT 415.120000 436.660000 416.320000 437.140000 ;
        RECT 415.120000 431.220000 416.320000 431.700000 ;
        RECT 460.120000 414.900000 461.320000 415.380000 ;
        RECT 460.120000 420.340000 461.320000 420.820000 ;
        RECT 460.120000 425.780000 461.320000 426.260000 ;
        RECT 460.120000 442.100000 461.320000 442.580000 ;
        RECT 460.120000 436.660000 461.320000 437.140000 ;
        RECT 460.120000 431.220000 461.320000 431.700000 ;
        RECT 415.120000 463.860000 416.320000 464.340000 ;
        RECT 415.120000 447.540000 416.320000 448.020000 ;
        RECT 415.120000 452.980000 416.320000 453.460000 ;
        RECT 415.120000 458.420000 416.320000 458.900000 ;
        RECT 415.120000 480.180000 416.320000 480.660000 ;
        RECT 415.120000 474.740000 416.320000 475.220000 ;
        RECT 415.120000 469.300000 416.320000 469.780000 ;
        RECT 460.120000 463.860000 461.320000 464.340000 ;
        RECT 460.120000 447.540000 461.320000 448.020000 ;
        RECT 460.120000 452.980000 461.320000 453.460000 ;
        RECT 460.120000 458.420000 461.320000 458.900000 ;
        RECT 460.120000 480.180000 461.320000 480.660000 ;
        RECT 460.120000 474.740000 461.320000 475.220000 ;
        RECT 460.120000 469.300000 461.320000 469.780000 ;
        RECT 505.120000 425.780000 506.320000 426.260000 ;
        RECT 505.120000 420.340000 506.320000 420.820000 ;
        RECT 505.120000 414.900000 506.320000 415.380000 ;
        RECT 505.120000 442.100000 506.320000 442.580000 ;
        RECT 505.120000 431.220000 506.320000 431.700000 ;
        RECT 505.120000 436.660000 506.320000 437.140000 ;
        RECT 545.600000 425.780000 546.800000 426.260000 ;
        RECT 545.600000 414.900000 546.800000 415.380000 ;
        RECT 545.600000 420.340000 546.800000 420.820000 ;
        RECT 545.600000 442.100000 546.800000 442.580000 ;
        RECT 545.600000 436.660000 546.800000 437.140000 ;
        RECT 545.600000 431.220000 546.800000 431.700000 ;
        RECT 505.120000 463.860000 506.320000 464.340000 ;
        RECT 505.120000 458.420000 506.320000 458.900000 ;
        RECT 505.120000 452.980000 506.320000 453.460000 ;
        RECT 505.120000 447.540000 506.320000 448.020000 ;
        RECT 505.120000 480.180000 506.320000 480.660000 ;
        RECT 505.120000 474.740000 506.320000 475.220000 ;
        RECT 505.120000 469.300000 506.320000 469.780000 ;
        RECT 545.600000 463.860000 546.800000 464.340000 ;
        RECT 545.600000 458.420000 546.800000 458.900000 ;
        RECT 545.600000 447.540000 546.800000 448.020000 ;
        RECT 545.600000 452.980000 546.800000 453.460000 ;
        RECT 545.600000 480.180000 546.800000 480.660000 ;
        RECT 545.600000 474.740000 546.800000 475.220000 ;
        RECT 545.600000 469.300000 546.800000 469.780000 ;
        RECT 415.120000 485.620000 416.320000 486.100000 ;
        RECT 415.120000 491.060000 416.320000 491.540000 ;
        RECT 415.120000 496.500000 416.320000 496.980000 ;
        RECT 415.120000 512.820000 416.320000 513.300000 ;
        RECT 415.120000 507.380000 416.320000 507.860000 ;
        RECT 415.120000 501.940000 416.320000 502.420000 ;
        RECT 460.120000 485.620000 461.320000 486.100000 ;
        RECT 460.120000 491.060000 461.320000 491.540000 ;
        RECT 460.120000 496.500000 461.320000 496.980000 ;
        RECT 460.120000 512.820000 461.320000 513.300000 ;
        RECT 460.120000 507.380000 461.320000 507.860000 ;
        RECT 460.120000 501.940000 461.320000 502.420000 ;
        RECT 415.120000 534.580000 416.320000 535.060000 ;
        RECT 415.120000 529.140000 416.320000 529.620000 ;
        RECT 415.120000 523.700000 416.320000 524.180000 ;
        RECT 415.120000 518.260000 416.320000 518.740000 ;
        RECT 460.120000 534.580000 461.320000 535.060000 ;
        RECT 460.120000 529.140000 461.320000 529.620000 ;
        RECT 460.120000 523.700000 461.320000 524.180000 ;
        RECT 460.120000 518.260000 461.320000 518.740000 ;
        RECT 505.120000 496.500000 506.320000 496.980000 ;
        RECT 505.120000 491.060000 506.320000 491.540000 ;
        RECT 505.120000 485.620000 506.320000 486.100000 ;
        RECT 505.120000 512.820000 506.320000 513.300000 ;
        RECT 505.120000 501.940000 506.320000 502.420000 ;
        RECT 505.120000 507.380000 506.320000 507.860000 ;
        RECT 545.600000 496.500000 546.800000 496.980000 ;
        RECT 545.600000 485.620000 546.800000 486.100000 ;
        RECT 545.600000 491.060000 546.800000 491.540000 ;
        RECT 545.600000 512.820000 546.800000 513.300000 ;
        RECT 545.600000 507.380000 546.800000 507.860000 ;
        RECT 545.600000 501.940000 546.800000 502.420000 ;
        RECT 505.120000 518.260000 506.320000 518.740000 ;
        RECT 505.120000 523.700000 506.320000 524.180000 ;
        RECT 505.120000 529.140000 506.320000 529.620000 ;
        RECT 505.120000 534.580000 506.320000 535.060000 ;
        RECT 545.600000 518.260000 546.800000 518.740000 ;
        RECT 545.600000 523.700000 546.800000 524.180000 ;
        RECT 545.600000 529.140000 546.800000 529.620000 ;
        RECT 545.600000 534.580000 546.800000 535.060000 ;
      LAYER met4 ;
        RECT 505.120000 3.230000 506.320000 545.360000 ;
        RECT 460.120000 3.230000 461.320000 545.360000 ;
        RECT 415.120000 3.230000 416.320000 545.360000 ;
        RECT 370.120000 3.230000 371.320000 545.360000 ;
        RECT 325.120000 3.230000 326.320000 545.360000 ;
        RECT 280.120000 3.230000 281.320000 545.360000 ;
        RECT 235.120000 3.230000 236.320000 545.360000 ;
        RECT 190.120000 3.230000 191.320000 545.360000 ;
        RECT 145.120000 3.230000 146.320000 545.360000 ;
        RECT 100.120000 3.230000 101.320000 545.360000 ;
        RECT 55.120000 3.230000 56.320000 545.360000 ;
        RECT 10.120000 3.230000 11.320000 545.360000 ;
        RECT 545.600000 0.000000 546.800000 549.780000 ;
        RECT 3.360000 0.000000 4.560000 549.780000 ;
        RECT 9.955000 34.100000 11.320000 34.580000 ;
        RECT 9.955000 12.340000 11.320000 12.820000 ;
        RECT 9.955000 23.220000 11.320000 23.700000 ;
        RECT 9.955000 17.780000 11.320000 18.260000 ;
        RECT 9.955000 28.660000 11.320000 29.140000 ;
        RECT 9.955000 39.540000 11.320000 40.020000 ;
        RECT 9.955000 50.420000 11.320000 50.900000 ;
        RECT 9.955000 44.980000 11.320000 45.460000 ;
        RECT 9.955000 55.860000 11.320000 56.340000 ;
        RECT 9.955000 66.740000 11.320000 67.220000 ;
        RECT 9.955000 61.300000 11.320000 61.780000 ;
        RECT 9.955000 72.180000 11.320000 72.660000 ;
        RECT 9.955000 83.060000 11.320000 83.540000 ;
        RECT 9.955000 77.620000 11.320000 78.100000 ;
        RECT 9.955000 93.940000 11.320000 94.420000 ;
        RECT 9.955000 88.500000 11.320000 88.980000 ;
        RECT 9.955000 99.380000 11.320000 99.860000 ;
        RECT 9.955000 110.260000 11.320000 110.740000 ;
        RECT 9.955000 104.820000 11.320000 105.300000 ;
        RECT 9.955000 115.700000 11.320000 116.180000 ;
        RECT 9.955000 126.580000 11.320000 127.060000 ;
        RECT 9.955000 121.140000 11.320000 121.620000 ;
        RECT 9.955000 132.020000 11.320000 132.500000 ;
        RECT 9.955000 142.900000 11.320000 143.380000 ;
        RECT 9.955000 137.460000 11.320000 137.940000 ;
        RECT 9.955000 153.780000 11.320000 154.260000 ;
        RECT 9.955000 148.340000 11.320000 148.820000 ;
        RECT 9.955000 159.220000 11.320000 159.700000 ;
        RECT 9.955000 170.100000 11.320000 170.580000 ;
        RECT 9.955000 164.660000 11.320000 165.140000 ;
        RECT 9.955000 175.540000 11.320000 176.020000 ;
        RECT 9.955000 186.420000 11.320000 186.900000 ;
        RECT 9.955000 180.980000 11.320000 181.460000 ;
        RECT 9.955000 197.300000 11.320000 197.780000 ;
        RECT 9.955000 191.860000 11.320000 192.340000 ;
        RECT 9.955000 202.740000 11.320000 203.220000 ;
        RECT 9.955000 213.620000 11.320000 214.100000 ;
        RECT 9.955000 208.180000 11.320000 208.660000 ;
        RECT 9.955000 219.060000 11.320000 219.540000 ;
        RECT 9.955000 229.940000 11.320000 230.420000 ;
        RECT 9.955000 224.500000 11.320000 224.980000 ;
        RECT 9.955000 235.380000 11.320000 235.860000 ;
        RECT 9.955000 246.260000 11.320000 246.740000 ;
        RECT 9.955000 240.820000 11.320000 241.300000 ;
        RECT 9.955000 257.140000 11.320000 257.620000 ;
        RECT 9.955000 251.700000 11.320000 252.180000 ;
        RECT 9.955000 262.580000 11.320000 263.060000 ;
        RECT 9.955000 273.460000 11.320000 273.940000 ;
        RECT 9.955000 268.020000 11.320000 268.500000 ;
        RECT 9.955000 278.900000 11.320000 279.380000 ;
        RECT 9.955000 289.780000 11.320000 290.260000 ;
        RECT 9.955000 284.340000 11.320000 284.820000 ;
        RECT 9.955000 300.660000 11.320000 301.140000 ;
        RECT 9.955000 295.220000 11.320000 295.700000 ;
        RECT 9.955000 306.100000 11.320000 306.580000 ;
        RECT 9.955000 316.980000 11.320000 317.460000 ;
        RECT 9.955000 311.540000 11.320000 312.020000 ;
        RECT 9.955000 322.420000 11.320000 322.900000 ;
        RECT 9.955000 333.300000 11.320000 333.780000 ;
        RECT 9.955000 327.860000 11.320000 328.340000 ;
        RECT 9.955000 338.740000 11.320000 339.220000 ;
        RECT 9.955000 360.500000 11.320000 360.980000 ;
        RECT 9.955000 349.620000 11.320000 350.100000 ;
        RECT 9.955000 344.180000 11.320000 344.660000 ;
        RECT 9.955000 355.060000 11.320000 355.540000 ;
        RECT 9.955000 365.940000 11.320000 366.420000 ;
        RECT 9.955000 376.820000 11.320000 377.300000 ;
        RECT 9.955000 371.380000 11.320000 371.860000 ;
        RECT 9.955000 382.260000 11.320000 382.740000 ;
        RECT 9.955000 393.140000 11.320000 393.620000 ;
        RECT 9.955000 387.700000 11.320000 388.180000 ;
        RECT 9.955000 398.580000 11.320000 399.060000 ;
        RECT 9.955000 409.460000 11.320000 409.940000 ;
        RECT 9.955000 404.020000 11.320000 404.500000 ;
        RECT 9.955000 420.340000 11.320000 420.820000 ;
        RECT 9.955000 414.900000 11.320000 415.380000 ;
        RECT 9.955000 425.780000 11.320000 426.260000 ;
        RECT 9.955000 436.660000 11.320000 437.140000 ;
        RECT 9.955000 431.220000 11.320000 431.700000 ;
        RECT 9.955000 442.100000 11.320000 442.580000 ;
        RECT 9.955000 463.860000 11.320000 464.340000 ;
        RECT 9.955000 452.980000 11.320000 453.460000 ;
        RECT 9.955000 447.540000 11.320000 448.020000 ;
        RECT 9.955000 458.420000 11.320000 458.900000 ;
        RECT 9.955000 469.300000 11.320000 469.780000 ;
        RECT 9.955000 480.180000 11.320000 480.660000 ;
        RECT 9.955000 474.740000 11.320000 475.220000 ;
        RECT 9.955000 485.620000 11.320000 486.100000 ;
        RECT 9.955000 496.500000 11.320000 496.980000 ;
        RECT 9.955000 491.060000 11.320000 491.540000 ;
        RECT 9.955000 501.940000 11.320000 502.420000 ;
        RECT 9.955000 512.820000 11.320000 513.300000 ;
        RECT 9.955000 507.380000 11.320000 507.860000 ;
        RECT 9.955000 523.700000 11.320000 524.180000 ;
        RECT 9.955000 518.260000 11.320000 518.740000 ;
        RECT 9.955000 529.140000 11.320000 529.620000 ;
        RECT 9.955000 534.580000 11.320000 535.060000 ;
    END
# end of P/G power stripe data as pin

  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 550.160000 549.780000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 550.160000 549.780000 ;
    LAYER met2 ;
      RECT 0.000000 1.040000 550.160000 549.780000 ;
      RECT 539.680000 0.000000 550.160000 1.040000 ;
      RECT 537.840000 0.000000 539.020000 1.040000 ;
      RECT 535.540000 0.000000 537.180000 1.040000 ;
      RECT 533.240000 0.000000 534.880000 1.040000 ;
      RECT 530.940000 0.000000 532.580000 1.040000 ;
      RECT 528.640000 0.000000 530.280000 1.040000 ;
      RECT 526.340000 0.000000 527.980000 1.040000 ;
      RECT 524.040000 0.000000 525.680000 1.040000 ;
      RECT 521.740000 0.000000 523.380000 1.040000 ;
      RECT 519.440000 0.000000 521.080000 1.040000 ;
      RECT 517.140000 0.000000 518.780000 1.040000 ;
      RECT 514.840000 0.000000 516.480000 1.040000 ;
      RECT 512.540000 0.000000 514.180000 1.040000 ;
      RECT 510.240000 0.000000 511.880000 1.040000 ;
      RECT 507.940000 0.000000 509.580000 1.040000 ;
      RECT 505.640000 0.000000 507.280000 1.040000 ;
      RECT 503.340000 0.000000 504.980000 1.040000 ;
      RECT 501.040000 0.000000 502.680000 1.040000 ;
      RECT 498.740000 0.000000 500.380000 1.040000 ;
      RECT 496.440000 0.000000 498.080000 1.040000 ;
      RECT 494.140000 0.000000 495.780000 1.040000 ;
      RECT 491.840000 0.000000 493.480000 1.040000 ;
      RECT 489.540000 0.000000 491.180000 1.040000 ;
      RECT 487.240000 0.000000 488.880000 1.040000 ;
      RECT 484.940000 0.000000 486.580000 1.040000 ;
      RECT 482.640000 0.000000 484.280000 1.040000 ;
      RECT 480.340000 0.000000 481.980000 1.040000 ;
      RECT 478.040000 0.000000 479.680000 1.040000 ;
      RECT 475.740000 0.000000 477.380000 1.040000 ;
      RECT 473.440000 0.000000 475.080000 1.040000 ;
      RECT 471.140000 0.000000 472.780000 1.040000 ;
      RECT 468.840000 0.000000 470.480000 1.040000 ;
      RECT 466.540000 0.000000 468.180000 1.040000 ;
      RECT 464.240000 0.000000 465.880000 1.040000 ;
      RECT 461.940000 0.000000 463.580000 1.040000 ;
      RECT 459.640000 0.000000 461.280000 1.040000 ;
      RECT 457.340000 0.000000 458.980000 1.040000 ;
      RECT 455.040000 0.000000 456.680000 1.040000 ;
      RECT 452.740000 0.000000 454.380000 1.040000 ;
      RECT 450.440000 0.000000 452.080000 1.040000 ;
      RECT 448.140000 0.000000 449.780000 1.040000 ;
      RECT 445.840000 0.000000 447.480000 1.040000 ;
      RECT 443.540000 0.000000 445.180000 1.040000 ;
      RECT 441.240000 0.000000 442.880000 1.040000 ;
      RECT 438.940000 0.000000 440.580000 1.040000 ;
      RECT 436.640000 0.000000 438.280000 1.040000 ;
      RECT 434.340000 0.000000 435.980000 1.040000 ;
      RECT 432.040000 0.000000 433.680000 1.040000 ;
      RECT 429.740000 0.000000 431.380000 1.040000 ;
      RECT 427.440000 0.000000 429.080000 1.040000 ;
      RECT 425.140000 0.000000 426.780000 1.040000 ;
      RECT 422.840000 0.000000 424.480000 1.040000 ;
      RECT 420.540000 0.000000 422.180000 1.040000 ;
      RECT 418.240000 0.000000 419.880000 1.040000 ;
      RECT 415.940000 0.000000 417.580000 1.040000 ;
      RECT 413.640000 0.000000 415.280000 1.040000 ;
      RECT 411.340000 0.000000 412.980000 1.040000 ;
      RECT 409.040000 0.000000 410.680000 1.040000 ;
      RECT 407.200000 0.000000 408.380000 1.040000 ;
      RECT 404.900000 0.000000 406.540000 1.040000 ;
      RECT 402.600000 0.000000 404.240000 1.040000 ;
      RECT 400.300000 0.000000 401.940000 1.040000 ;
      RECT 398.000000 0.000000 399.640000 1.040000 ;
      RECT 395.700000 0.000000 397.340000 1.040000 ;
      RECT 393.400000 0.000000 395.040000 1.040000 ;
      RECT 391.100000 0.000000 392.740000 1.040000 ;
      RECT 388.800000 0.000000 390.440000 1.040000 ;
      RECT 386.500000 0.000000 388.140000 1.040000 ;
      RECT 384.200000 0.000000 385.840000 1.040000 ;
      RECT 381.900000 0.000000 383.540000 1.040000 ;
      RECT 379.600000 0.000000 381.240000 1.040000 ;
      RECT 377.300000 0.000000 378.940000 1.040000 ;
      RECT 375.000000 0.000000 376.640000 1.040000 ;
      RECT 372.700000 0.000000 374.340000 1.040000 ;
      RECT 370.400000 0.000000 372.040000 1.040000 ;
      RECT 368.100000 0.000000 369.740000 1.040000 ;
      RECT 365.800000 0.000000 367.440000 1.040000 ;
      RECT 363.500000 0.000000 365.140000 1.040000 ;
      RECT 361.200000 0.000000 362.840000 1.040000 ;
      RECT 358.900000 0.000000 360.540000 1.040000 ;
      RECT 356.600000 0.000000 358.240000 1.040000 ;
      RECT 354.300000 0.000000 355.940000 1.040000 ;
      RECT 352.000000 0.000000 353.640000 1.040000 ;
      RECT 349.700000 0.000000 351.340000 1.040000 ;
      RECT 347.400000 0.000000 349.040000 1.040000 ;
      RECT 345.100000 0.000000 346.740000 1.040000 ;
      RECT 342.800000 0.000000 344.440000 1.040000 ;
      RECT 340.500000 0.000000 342.140000 1.040000 ;
      RECT 338.200000 0.000000 339.840000 1.040000 ;
      RECT 335.900000 0.000000 337.540000 1.040000 ;
      RECT 333.600000 0.000000 335.240000 1.040000 ;
      RECT 331.300000 0.000000 332.940000 1.040000 ;
      RECT 329.000000 0.000000 330.640000 1.040000 ;
      RECT 326.700000 0.000000 328.340000 1.040000 ;
      RECT 324.400000 0.000000 326.040000 1.040000 ;
      RECT 322.100000 0.000000 323.740000 1.040000 ;
      RECT 319.800000 0.000000 321.440000 1.040000 ;
      RECT 317.500000 0.000000 319.140000 1.040000 ;
      RECT 315.200000 0.000000 316.840000 1.040000 ;
      RECT 312.900000 0.000000 314.540000 1.040000 ;
      RECT 310.600000 0.000000 312.240000 1.040000 ;
      RECT 308.300000 0.000000 309.940000 1.040000 ;
      RECT 306.000000 0.000000 307.640000 1.040000 ;
      RECT 303.700000 0.000000 305.340000 1.040000 ;
      RECT 301.400000 0.000000 303.040000 1.040000 ;
      RECT 299.100000 0.000000 300.740000 1.040000 ;
      RECT 296.800000 0.000000 298.440000 1.040000 ;
      RECT 294.500000 0.000000 296.140000 1.040000 ;
      RECT 292.200000 0.000000 293.840000 1.040000 ;
      RECT 289.900000 0.000000 291.540000 1.040000 ;
      RECT 287.600000 0.000000 289.240000 1.040000 ;
      RECT 285.300000 0.000000 286.940000 1.040000 ;
      RECT 283.000000 0.000000 284.640000 1.040000 ;
      RECT 280.700000 0.000000 282.340000 1.040000 ;
      RECT 278.400000 0.000000 280.040000 1.040000 ;
      RECT 276.100000 0.000000 277.740000 1.040000 ;
      RECT 274.260000 0.000000 275.440000 1.040000 ;
      RECT 271.960000 0.000000 273.600000 1.040000 ;
      RECT 269.660000 0.000000 271.300000 1.040000 ;
      RECT 267.360000 0.000000 269.000000 1.040000 ;
      RECT 265.060000 0.000000 266.700000 1.040000 ;
      RECT 262.760000 0.000000 264.400000 1.040000 ;
      RECT 260.460000 0.000000 262.100000 1.040000 ;
      RECT 258.160000 0.000000 259.800000 1.040000 ;
      RECT 255.860000 0.000000 257.500000 1.040000 ;
      RECT 253.560000 0.000000 255.200000 1.040000 ;
      RECT 251.260000 0.000000 252.900000 1.040000 ;
      RECT 248.960000 0.000000 250.600000 1.040000 ;
      RECT 246.660000 0.000000 248.300000 1.040000 ;
      RECT 244.360000 0.000000 246.000000 1.040000 ;
      RECT 242.060000 0.000000 243.700000 1.040000 ;
      RECT 239.760000 0.000000 241.400000 1.040000 ;
      RECT 237.460000 0.000000 239.100000 1.040000 ;
      RECT 235.160000 0.000000 236.800000 1.040000 ;
      RECT 232.860000 0.000000 234.500000 1.040000 ;
      RECT 230.560000 0.000000 232.200000 1.040000 ;
      RECT 228.260000 0.000000 229.900000 1.040000 ;
      RECT 225.960000 0.000000 227.600000 1.040000 ;
      RECT 223.660000 0.000000 225.300000 1.040000 ;
      RECT 221.360000 0.000000 223.000000 1.040000 ;
      RECT 219.060000 0.000000 220.700000 1.040000 ;
      RECT 216.760000 0.000000 218.400000 1.040000 ;
      RECT 214.460000 0.000000 216.100000 1.040000 ;
      RECT 212.160000 0.000000 213.800000 1.040000 ;
      RECT 209.860000 0.000000 211.500000 1.040000 ;
      RECT 207.560000 0.000000 209.200000 1.040000 ;
      RECT 205.260000 0.000000 206.900000 1.040000 ;
      RECT 202.960000 0.000000 204.600000 1.040000 ;
      RECT 200.660000 0.000000 202.300000 1.040000 ;
      RECT 198.360000 0.000000 200.000000 1.040000 ;
      RECT 196.060000 0.000000 197.700000 1.040000 ;
      RECT 193.760000 0.000000 195.400000 1.040000 ;
      RECT 191.460000 0.000000 193.100000 1.040000 ;
      RECT 189.160000 0.000000 190.800000 1.040000 ;
      RECT 186.860000 0.000000 188.500000 1.040000 ;
      RECT 184.560000 0.000000 186.200000 1.040000 ;
      RECT 182.260000 0.000000 183.900000 1.040000 ;
      RECT 179.960000 0.000000 181.600000 1.040000 ;
      RECT 177.660000 0.000000 179.300000 1.040000 ;
      RECT 175.360000 0.000000 177.000000 1.040000 ;
      RECT 173.060000 0.000000 174.700000 1.040000 ;
      RECT 170.760000 0.000000 172.400000 1.040000 ;
      RECT 168.460000 0.000000 170.100000 1.040000 ;
      RECT 166.160000 0.000000 167.800000 1.040000 ;
      RECT 163.860000 0.000000 165.500000 1.040000 ;
      RECT 161.560000 0.000000 163.200000 1.040000 ;
      RECT 159.260000 0.000000 160.900000 1.040000 ;
      RECT 156.960000 0.000000 158.600000 1.040000 ;
      RECT 154.660000 0.000000 156.300000 1.040000 ;
      RECT 152.360000 0.000000 154.000000 1.040000 ;
      RECT 150.060000 0.000000 151.700000 1.040000 ;
      RECT 147.760000 0.000000 149.400000 1.040000 ;
      RECT 145.460000 0.000000 147.100000 1.040000 ;
      RECT 143.160000 0.000000 144.800000 1.040000 ;
      RECT 141.320000 0.000000 142.500000 1.040000 ;
      RECT 139.020000 0.000000 140.660000 1.040000 ;
      RECT 136.720000 0.000000 138.360000 1.040000 ;
      RECT 134.420000 0.000000 136.060000 1.040000 ;
      RECT 132.120000 0.000000 133.760000 1.040000 ;
      RECT 129.820000 0.000000 131.460000 1.040000 ;
      RECT 127.520000 0.000000 129.160000 1.040000 ;
      RECT 125.220000 0.000000 126.860000 1.040000 ;
      RECT 122.920000 0.000000 124.560000 1.040000 ;
      RECT 120.620000 0.000000 122.260000 1.040000 ;
      RECT 118.320000 0.000000 119.960000 1.040000 ;
      RECT 116.020000 0.000000 117.660000 1.040000 ;
      RECT 113.720000 0.000000 115.360000 1.040000 ;
      RECT 111.420000 0.000000 113.060000 1.040000 ;
      RECT 109.120000 0.000000 110.760000 1.040000 ;
      RECT 106.820000 0.000000 108.460000 1.040000 ;
      RECT 104.520000 0.000000 106.160000 1.040000 ;
      RECT 102.220000 0.000000 103.860000 1.040000 ;
      RECT 99.920000 0.000000 101.560000 1.040000 ;
      RECT 97.620000 0.000000 99.260000 1.040000 ;
      RECT 95.320000 0.000000 96.960000 1.040000 ;
      RECT 93.020000 0.000000 94.660000 1.040000 ;
      RECT 90.720000 0.000000 92.360000 1.040000 ;
      RECT 88.420000 0.000000 90.060000 1.040000 ;
      RECT 86.120000 0.000000 87.760000 1.040000 ;
      RECT 83.820000 0.000000 85.460000 1.040000 ;
      RECT 81.520000 0.000000 83.160000 1.040000 ;
      RECT 79.220000 0.000000 80.860000 1.040000 ;
      RECT 76.920000 0.000000 78.560000 1.040000 ;
      RECT 74.620000 0.000000 76.260000 1.040000 ;
      RECT 72.320000 0.000000 73.960000 1.040000 ;
      RECT 70.020000 0.000000 71.660000 1.040000 ;
      RECT 67.720000 0.000000 69.360000 1.040000 ;
      RECT 65.420000 0.000000 67.060000 1.040000 ;
      RECT 63.120000 0.000000 64.760000 1.040000 ;
      RECT 60.820000 0.000000 62.460000 1.040000 ;
      RECT 58.520000 0.000000 60.160000 1.040000 ;
      RECT 56.220000 0.000000 57.860000 1.040000 ;
      RECT 53.920000 0.000000 55.560000 1.040000 ;
      RECT 51.620000 0.000000 53.260000 1.040000 ;
      RECT 49.320000 0.000000 50.960000 1.040000 ;
      RECT 47.020000 0.000000 48.660000 1.040000 ;
      RECT 44.720000 0.000000 46.360000 1.040000 ;
      RECT 42.420000 0.000000 44.060000 1.040000 ;
      RECT 40.120000 0.000000 41.760000 1.040000 ;
      RECT 37.820000 0.000000 39.460000 1.040000 ;
      RECT 35.520000 0.000000 37.160000 1.040000 ;
      RECT 33.220000 0.000000 34.860000 1.040000 ;
      RECT 30.920000 0.000000 32.560000 1.040000 ;
      RECT 28.620000 0.000000 30.260000 1.040000 ;
      RECT 26.320000 0.000000 27.960000 1.040000 ;
      RECT 24.020000 0.000000 25.660000 1.040000 ;
      RECT 21.720000 0.000000 23.360000 1.040000 ;
      RECT 19.420000 0.000000 21.060000 1.040000 ;
      RECT 17.120000 0.000000 18.760000 1.040000 ;
      RECT 14.820000 0.000000 16.460000 1.040000 ;
      RECT 12.520000 0.000000 14.160000 1.040000 ;
      RECT 10.680000 0.000000 11.860000 1.040000 ;
      RECT 0.000000 0.000000 10.020000 1.040000 ;
    LAYER met3 ;
      RECT 0.000000 545.660000 550.160000 549.780000 ;
      RECT 0.000000 543.460000 550.160000 543.860000 ;
      RECT 0.000000 539.390000 550.160000 541.660000 ;
      RECT 0.000000 538.410000 548.960000 539.390000 ;
      RECT 0.000000 538.080000 550.160000 538.410000 ;
      RECT 544.900000 537.000000 550.160000 538.080000 ;
      RECT 508.620000 537.000000 543.100000 538.080000 ;
      RECT 463.620000 537.000000 506.820000 538.080000 ;
      RECT 418.620000 537.000000 461.820000 538.080000 ;
      RECT 373.620000 537.000000 416.820000 538.080000 ;
      RECT 328.620000 537.000000 371.820000 538.080000 ;
      RECT 283.620000 537.000000 326.820000 538.080000 ;
      RECT 238.620000 537.000000 281.820000 538.080000 ;
      RECT 193.620000 537.000000 236.820000 538.080000 ;
      RECT 148.620000 537.000000 191.820000 538.080000 ;
      RECT 103.620000 537.000000 146.820000 538.080000 ;
      RECT 58.620000 537.000000 101.820000 538.080000 ;
      RECT 13.620000 537.000000 56.820000 538.080000 ;
      RECT 7.060000 537.000000 11.820000 538.080000 ;
      RECT 0.000000 537.000000 5.260000 538.080000 ;
      RECT 0.000000 536.340000 550.160000 537.000000 ;
      RECT 0.000000 535.360000 548.960000 536.340000 ;
      RECT 547.100000 534.280000 550.160000 535.360000 ;
      RECT 506.620000 534.280000 545.300000 535.360000 ;
      RECT 461.620000 534.280000 504.820000 535.360000 ;
      RECT 416.620000 534.280000 459.820000 535.360000 ;
      RECT 371.620000 534.280000 414.820000 535.360000 ;
      RECT 326.620000 534.280000 369.820000 535.360000 ;
      RECT 281.620000 534.280000 324.820000 535.360000 ;
      RECT 236.620000 534.280000 279.820000 535.360000 ;
      RECT 191.620000 534.280000 234.820000 535.360000 ;
      RECT 146.620000 534.280000 189.820000 535.360000 ;
      RECT 101.620000 534.280000 144.820000 535.360000 ;
      RECT 56.620000 534.280000 99.820000 535.360000 ;
      RECT 11.620000 534.280000 54.820000 535.360000 ;
      RECT 4.860000 534.280000 9.655000 535.360000 ;
      RECT 0.000000 534.280000 3.060000 535.360000 ;
      RECT 0.000000 533.290000 550.160000 534.280000 ;
      RECT 0.000000 532.640000 548.960000 533.290000 ;
      RECT 544.900000 532.310000 548.960000 532.640000 ;
      RECT 544.900000 531.560000 550.160000 532.310000 ;
      RECT 508.620000 531.560000 543.100000 532.640000 ;
      RECT 463.620000 531.560000 506.820000 532.640000 ;
      RECT 418.620000 531.560000 461.820000 532.640000 ;
      RECT 373.620000 531.560000 416.820000 532.640000 ;
      RECT 328.620000 531.560000 371.820000 532.640000 ;
      RECT 283.620000 531.560000 326.820000 532.640000 ;
      RECT 238.620000 531.560000 281.820000 532.640000 ;
      RECT 193.620000 531.560000 236.820000 532.640000 ;
      RECT 148.620000 531.560000 191.820000 532.640000 ;
      RECT 103.620000 531.560000 146.820000 532.640000 ;
      RECT 58.620000 531.560000 101.820000 532.640000 ;
      RECT 13.620000 531.560000 56.820000 532.640000 ;
      RECT 7.060000 531.560000 11.820000 532.640000 ;
      RECT 0.000000 531.560000 5.260000 532.640000 ;
      RECT 0.000000 530.240000 550.160000 531.560000 ;
      RECT 0.000000 529.920000 548.960000 530.240000 ;
      RECT 547.100000 529.260000 548.960000 529.920000 ;
      RECT 547.100000 528.840000 550.160000 529.260000 ;
      RECT 506.620000 528.840000 545.300000 529.920000 ;
      RECT 461.620000 528.840000 504.820000 529.920000 ;
      RECT 416.620000 528.840000 459.820000 529.920000 ;
      RECT 371.620000 528.840000 414.820000 529.920000 ;
      RECT 326.620000 528.840000 369.820000 529.920000 ;
      RECT 281.620000 528.840000 324.820000 529.920000 ;
      RECT 236.620000 528.840000 279.820000 529.920000 ;
      RECT 191.620000 528.840000 234.820000 529.920000 ;
      RECT 146.620000 528.840000 189.820000 529.920000 ;
      RECT 101.620000 528.840000 144.820000 529.920000 ;
      RECT 56.620000 528.840000 99.820000 529.920000 ;
      RECT 11.620000 528.840000 54.820000 529.920000 ;
      RECT 4.860000 528.840000 9.655000 529.920000 ;
      RECT 0.000000 528.840000 3.060000 529.920000 ;
      RECT 0.000000 527.200000 550.160000 528.840000 ;
      RECT 544.900000 527.190000 550.160000 527.200000 ;
      RECT 544.900000 526.210000 548.960000 527.190000 ;
      RECT 544.900000 526.120000 550.160000 526.210000 ;
      RECT 508.620000 526.120000 543.100000 527.200000 ;
      RECT 463.620000 526.120000 506.820000 527.200000 ;
      RECT 418.620000 526.120000 461.820000 527.200000 ;
      RECT 373.620000 526.120000 416.820000 527.200000 ;
      RECT 328.620000 526.120000 371.820000 527.200000 ;
      RECT 283.620000 526.120000 326.820000 527.200000 ;
      RECT 238.620000 526.120000 281.820000 527.200000 ;
      RECT 193.620000 526.120000 236.820000 527.200000 ;
      RECT 148.620000 526.120000 191.820000 527.200000 ;
      RECT 103.620000 526.120000 146.820000 527.200000 ;
      RECT 58.620000 526.120000 101.820000 527.200000 ;
      RECT 13.620000 526.120000 56.820000 527.200000 ;
      RECT 7.060000 526.120000 11.820000 527.200000 ;
      RECT 0.000000 526.120000 5.260000 527.200000 ;
      RECT 0.000000 524.480000 550.160000 526.120000 ;
      RECT 547.100000 524.140000 550.160000 524.480000 ;
      RECT 547.100000 523.400000 548.960000 524.140000 ;
      RECT 506.620000 523.400000 545.300000 524.480000 ;
      RECT 461.620000 523.400000 504.820000 524.480000 ;
      RECT 416.620000 523.400000 459.820000 524.480000 ;
      RECT 371.620000 523.400000 414.820000 524.480000 ;
      RECT 326.620000 523.400000 369.820000 524.480000 ;
      RECT 281.620000 523.400000 324.820000 524.480000 ;
      RECT 236.620000 523.400000 279.820000 524.480000 ;
      RECT 191.620000 523.400000 234.820000 524.480000 ;
      RECT 146.620000 523.400000 189.820000 524.480000 ;
      RECT 101.620000 523.400000 144.820000 524.480000 ;
      RECT 56.620000 523.400000 99.820000 524.480000 ;
      RECT 11.620000 523.400000 54.820000 524.480000 ;
      RECT 4.860000 523.400000 9.655000 524.480000 ;
      RECT 0.000000 523.400000 3.060000 524.480000 ;
      RECT 0.000000 523.160000 548.960000 523.400000 ;
      RECT 0.000000 521.760000 550.160000 523.160000 ;
      RECT 544.900000 520.680000 550.160000 521.760000 ;
      RECT 508.620000 520.680000 543.100000 521.760000 ;
      RECT 463.620000 520.680000 506.820000 521.760000 ;
      RECT 418.620000 520.680000 461.820000 521.760000 ;
      RECT 373.620000 520.680000 416.820000 521.760000 ;
      RECT 328.620000 520.680000 371.820000 521.760000 ;
      RECT 283.620000 520.680000 326.820000 521.760000 ;
      RECT 238.620000 520.680000 281.820000 521.760000 ;
      RECT 193.620000 520.680000 236.820000 521.760000 ;
      RECT 148.620000 520.680000 191.820000 521.760000 ;
      RECT 103.620000 520.680000 146.820000 521.760000 ;
      RECT 58.620000 520.680000 101.820000 521.760000 ;
      RECT 13.620000 520.680000 56.820000 521.760000 ;
      RECT 7.060000 520.680000 11.820000 521.760000 ;
      RECT 0.000000 520.680000 5.260000 521.760000 ;
      RECT 0.000000 520.480000 550.160000 520.680000 ;
      RECT 0.000000 519.500000 548.960000 520.480000 ;
      RECT 0.000000 519.040000 550.160000 519.500000 ;
      RECT 547.100000 517.960000 550.160000 519.040000 ;
      RECT 506.620000 517.960000 545.300000 519.040000 ;
      RECT 461.620000 517.960000 504.820000 519.040000 ;
      RECT 416.620000 517.960000 459.820000 519.040000 ;
      RECT 371.620000 517.960000 414.820000 519.040000 ;
      RECT 326.620000 517.960000 369.820000 519.040000 ;
      RECT 281.620000 517.960000 324.820000 519.040000 ;
      RECT 236.620000 517.960000 279.820000 519.040000 ;
      RECT 191.620000 517.960000 234.820000 519.040000 ;
      RECT 146.620000 517.960000 189.820000 519.040000 ;
      RECT 101.620000 517.960000 144.820000 519.040000 ;
      RECT 56.620000 517.960000 99.820000 519.040000 ;
      RECT 11.620000 517.960000 54.820000 519.040000 ;
      RECT 4.860000 517.960000 9.655000 519.040000 ;
      RECT 0.000000 517.960000 3.060000 519.040000 ;
      RECT 0.000000 517.430000 550.160000 517.960000 ;
      RECT 0.000000 516.450000 548.960000 517.430000 ;
      RECT 0.000000 516.320000 550.160000 516.450000 ;
      RECT 544.900000 515.240000 550.160000 516.320000 ;
      RECT 508.620000 515.240000 543.100000 516.320000 ;
      RECT 463.620000 515.240000 506.820000 516.320000 ;
      RECT 418.620000 515.240000 461.820000 516.320000 ;
      RECT 373.620000 515.240000 416.820000 516.320000 ;
      RECT 328.620000 515.240000 371.820000 516.320000 ;
      RECT 283.620000 515.240000 326.820000 516.320000 ;
      RECT 238.620000 515.240000 281.820000 516.320000 ;
      RECT 193.620000 515.240000 236.820000 516.320000 ;
      RECT 148.620000 515.240000 191.820000 516.320000 ;
      RECT 103.620000 515.240000 146.820000 516.320000 ;
      RECT 58.620000 515.240000 101.820000 516.320000 ;
      RECT 13.620000 515.240000 56.820000 516.320000 ;
      RECT 7.060000 515.240000 11.820000 516.320000 ;
      RECT 0.000000 515.240000 5.260000 516.320000 ;
      RECT 0.000000 514.380000 550.160000 515.240000 ;
      RECT 0.000000 513.600000 548.960000 514.380000 ;
      RECT 547.100000 513.400000 548.960000 513.600000 ;
      RECT 547.100000 512.520000 550.160000 513.400000 ;
      RECT 506.620000 512.520000 545.300000 513.600000 ;
      RECT 461.620000 512.520000 504.820000 513.600000 ;
      RECT 416.620000 512.520000 459.820000 513.600000 ;
      RECT 371.620000 512.520000 414.820000 513.600000 ;
      RECT 326.620000 512.520000 369.820000 513.600000 ;
      RECT 281.620000 512.520000 324.820000 513.600000 ;
      RECT 236.620000 512.520000 279.820000 513.600000 ;
      RECT 191.620000 512.520000 234.820000 513.600000 ;
      RECT 146.620000 512.520000 189.820000 513.600000 ;
      RECT 101.620000 512.520000 144.820000 513.600000 ;
      RECT 56.620000 512.520000 99.820000 513.600000 ;
      RECT 11.620000 512.520000 54.820000 513.600000 ;
      RECT 4.860000 512.520000 9.655000 513.600000 ;
      RECT 0.000000 512.520000 3.060000 513.600000 ;
      RECT 0.000000 511.330000 550.160000 512.520000 ;
      RECT 0.000000 510.880000 548.960000 511.330000 ;
      RECT 544.900000 510.350000 548.960000 510.880000 ;
      RECT 544.900000 509.800000 550.160000 510.350000 ;
      RECT 508.620000 509.800000 543.100000 510.880000 ;
      RECT 463.620000 509.800000 506.820000 510.880000 ;
      RECT 418.620000 509.800000 461.820000 510.880000 ;
      RECT 373.620000 509.800000 416.820000 510.880000 ;
      RECT 328.620000 509.800000 371.820000 510.880000 ;
      RECT 283.620000 509.800000 326.820000 510.880000 ;
      RECT 238.620000 509.800000 281.820000 510.880000 ;
      RECT 193.620000 509.800000 236.820000 510.880000 ;
      RECT 148.620000 509.800000 191.820000 510.880000 ;
      RECT 103.620000 509.800000 146.820000 510.880000 ;
      RECT 58.620000 509.800000 101.820000 510.880000 ;
      RECT 13.620000 509.800000 56.820000 510.880000 ;
      RECT 7.060000 509.800000 11.820000 510.880000 ;
      RECT 0.000000 509.800000 5.260000 510.880000 ;
      RECT 0.000000 508.280000 550.160000 509.800000 ;
      RECT 0.000000 508.160000 548.960000 508.280000 ;
      RECT 547.100000 507.300000 548.960000 508.160000 ;
      RECT 547.100000 507.080000 550.160000 507.300000 ;
      RECT 506.620000 507.080000 545.300000 508.160000 ;
      RECT 461.620000 507.080000 504.820000 508.160000 ;
      RECT 416.620000 507.080000 459.820000 508.160000 ;
      RECT 371.620000 507.080000 414.820000 508.160000 ;
      RECT 326.620000 507.080000 369.820000 508.160000 ;
      RECT 281.620000 507.080000 324.820000 508.160000 ;
      RECT 236.620000 507.080000 279.820000 508.160000 ;
      RECT 191.620000 507.080000 234.820000 508.160000 ;
      RECT 146.620000 507.080000 189.820000 508.160000 ;
      RECT 101.620000 507.080000 144.820000 508.160000 ;
      RECT 56.620000 507.080000 99.820000 508.160000 ;
      RECT 11.620000 507.080000 54.820000 508.160000 ;
      RECT 4.860000 507.080000 9.655000 508.160000 ;
      RECT 0.000000 507.080000 3.060000 508.160000 ;
      RECT 0.000000 505.440000 550.160000 507.080000 ;
      RECT 544.900000 505.230000 550.160000 505.440000 ;
      RECT 544.900000 504.360000 548.960000 505.230000 ;
      RECT 508.620000 504.360000 543.100000 505.440000 ;
      RECT 463.620000 504.360000 506.820000 505.440000 ;
      RECT 418.620000 504.360000 461.820000 505.440000 ;
      RECT 373.620000 504.360000 416.820000 505.440000 ;
      RECT 328.620000 504.360000 371.820000 505.440000 ;
      RECT 283.620000 504.360000 326.820000 505.440000 ;
      RECT 238.620000 504.360000 281.820000 505.440000 ;
      RECT 193.620000 504.360000 236.820000 505.440000 ;
      RECT 148.620000 504.360000 191.820000 505.440000 ;
      RECT 103.620000 504.360000 146.820000 505.440000 ;
      RECT 58.620000 504.360000 101.820000 505.440000 ;
      RECT 13.620000 504.360000 56.820000 505.440000 ;
      RECT 7.060000 504.360000 11.820000 505.440000 ;
      RECT 0.000000 504.360000 5.260000 505.440000 ;
      RECT 0.000000 504.250000 548.960000 504.360000 ;
      RECT 0.000000 502.720000 550.160000 504.250000 ;
      RECT 547.100000 501.640000 550.160000 502.720000 ;
      RECT 506.620000 501.640000 545.300000 502.720000 ;
      RECT 461.620000 501.640000 504.820000 502.720000 ;
      RECT 416.620000 501.640000 459.820000 502.720000 ;
      RECT 371.620000 501.640000 414.820000 502.720000 ;
      RECT 326.620000 501.640000 369.820000 502.720000 ;
      RECT 281.620000 501.640000 324.820000 502.720000 ;
      RECT 236.620000 501.640000 279.820000 502.720000 ;
      RECT 191.620000 501.640000 234.820000 502.720000 ;
      RECT 146.620000 501.640000 189.820000 502.720000 ;
      RECT 101.620000 501.640000 144.820000 502.720000 ;
      RECT 56.620000 501.640000 99.820000 502.720000 ;
      RECT 11.620000 501.640000 54.820000 502.720000 ;
      RECT 4.860000 501.640000 9.655000 502.720000 ;
      RECT 0.000000 501.640000 3.060000 502.720000 ;
      RECT 0.000000 501.570000 550.160000 501.640000 ;
      RECT 0.000000 500.590000 548.960000 501.570000 ;
      RECT 0.000000 500.000000 550.160000 500.590000 ;
      RECT 544.900000 498.920000 550.160000 500.000000 ;
      RECT 508.620000 498.920000 543.100000 500.000000 ;
      RECT 463.620000 498.920000 506.820000 500.000000 ;
      RECT 418.620000 498.920000 461.820000 500.000000 ;
      RECT 373.620000 498.920000 416.820000 500.000000 ;
      RECT 328.620000 498.920000 371.820000 500.000000 ;
      RECT 283.620000 498.920000 326.820000 500.000000 ;
      RECT 238.620000 498.920000 281.820000 500.000000 ;
      RECT 193.620000 498.920000 236.820000 500.000000 ;
      RECT 148.620000 498.920000 191.820000 500.000000 ;
      RECT 103.620000 498.920000 146.820000 500.000000 ;
      RECT 58.620000 498.920000 101.820000 500.000000 ;
      RECT 13.620000 498.920000 56.820000 500.000000 ;
      RECT 7.060000 498.920000 11.820000 500.000000 ;
      RECT 0.000000 498.920000 5.260000 500.000000 ;
      RECT 0.000000 498.520000 550.160000 498.920000 ;
      RECT 0.000000 497.540000 548.960000 498.520000 ;
      RECT 0.000000 497.280000 550.160000 497.540000 ;
      RECT 547.100000 496.200000 550.160000 497.280000 ;
      RECT 506.620000 496.200000 545.300000 497.280000 ;
      RECT 461.620000 496.200000 504.820000 497.280000 ;
      RECT 416.620000 496.200000 459.820000 497.280000 ;
      RECT 371.620000 496.200000 414.820000 497.280000 ;
      RECT 326.620000 496.200000 369.820000 497.280000 ;
      RECT 281.620000 496.200000 324.820000 497.280000 ;
      RECT 236.620000 496.200000 279.820000 497.280000 ;
      RECT 191.620000 496.200000 234.820000 497.280000 ;
      RECT 146.620000 496.200000 189.820000 497.280000 ;
      RECT 101.620000 496.200000 144.820000 497.280000 ;
      RECT 56.620000 496.200000 99.820000 497.280000 ;
      RECT 11.620000 496.200000 54.820000 497.280000 ;
      RECT 4.860000 496.200000 9.655000 497.280000 ;
      RECT 0.000000 496.200000 3.060000 497.280000 ;
      RECT 0.000000 495.470000 550.160000 496.200000 ;
      RECT 0.000000 494.560000 548.960000 495.470000 ;
      RECT 544.900000 494.490000 548.960000 494.560000 ;
      RECT 544.900000 493.480000 550.160000 494.490000 ;
      RECT 508.620000 493.480000 543.100000 494.560000 ;
      RECT 463.620000 493.480000 506.820000 494.560000 ;
      RECT 418.620000 493.480000 461.820000 494.560000 ;
      RECT 373.620000 493.480000 416.820000 494.560000 ;
      RECT 328.620000 493.480000 371.820000 494.560000 ;
      RECT 283.620000 493.480000 326.820000 494.560000 ;
      RECT 238.620000 493.480000 281.820000 494.560000 ;
      RECT 193.620000 493.480000 236.820000 494.560000 ;
      RECT 148.620000 493.480000 191.820000 494.560000 ;
      RECT 103.620000 493.480000 146.820000 494.560000 ;
      RECT 58.620000 493.480000 101.820000 494.560000 ;
      RECT 13.620000 493.480000 56.820000 494.560000 ;
      RECT 7.060000 493.480000 11.820000 494.560000 ;
      RECT 0.000000 493.480000 5.260000 494.560000 ;
      RECT 0.000000 492.420000 550.160000 493.480000 ;
      RECT 0.000000 491.840000 548.960000 492.420000 ;
      RECT 547.100000 491.440000 548.960000 491.840000 ;
      RECT 547.100000 490.760000 550.160000 491.440000 ;
      RECT 506.620000 490.760000 545.300000 491.840000 ;
      RECT 461.620000 490.760000 504.820000 491.840000 ;
      RECT 416.620000 490.760000 459.820000 491.840000 ;
      RECT 371.620000 490.760000 414.820000 491.840000 ;
      RECT 326.620000 490.760000 369.820000 491.840000 ;
      RECT 281.620000 490.760000 324.820000 491.840000 ;
      RECT 236.620000 490.760000 279.820000 491.840000 ;
      RECT 191.620000 490.760000 234.820000 491.840000 ;
      RECT 146.620000 490.760000 189.820000 491.840000 ;
      RECT 101.620000 490.760000 144.820000 491.840000 ;
      RECT 56.620000 490.760000 99.820000 491.840000 ;
      RECT 11.620000 490.760000 54.820000 491.840000 ;
      RECT 4.860000 490.760000 9.655000 491.840000 ;
      RECT 0.000000 490.760000 3.060000 491.840000 ;
      RECT 0.000000 489.370000 550.160000 490.760000 ;
      RECT 0.000000 489.120000 548.960000 489.370000 ;
      RECT 544.900000 488.390000 548.960000 489.120000 ;
      RECT 544.900000 488.040000 550.160000 488.390000 ;
      RECT 508.620000 488.040000 543.100000 489.120000 ;
      RECT 463.620000 488.040000 506.820000 489.120000 ;
      RECT 418.620000 488.040000 461.820000 489.120000 ;
      RECT 373.620000 488.040000 416.820000 489.120000 ;
      RECT 328.620000 488.040000 371.820000 489.120000 ;
      RECT 283.620000 488.040000 326.820000 489.120000 ;
      RECT 238.620000 488.040000 281.820000 489.120000 ;
      RECT 193.620000 488.040000 236.820000 489.120000 ;
      RECT 148.620000 488.040000 191.820000 489.120000 ;
      RECT 103.620000 488.040000 146.820000 489.120000 ;
      RECT 58.620000 488.040000 101.820000 489.120000 ;
      RECT 13.620000 488.040000 56.820000 489.120000 ;
      RECT 7.060000 488.040000 11.820000 489.120000 ;
      RECT 0.000000 488.040000 5.260000 489.120000 ;
      RECT 0.000000 486.400000 550.160000 488.040000 ;
      RECT 547.100000 486.320000 550.160000 486.400000 ;
      RECT 547.100000 485.340000 548.960000 486.320000 ;
      RECT 547.100000 485.320000 550.160000 485.340000 ;
      RECT 506.620000 485.320000 545.300000 486.400000 ;
      RECT 461.620000 485.320000 504.820000 486.400000 ;
      RECT 416.620000 485.320000 459.820000 486.400000 ;
      RECT 371.620000 485.320000 414.820000 486.400000 ;
      RECT 326.620000 485.320000 369.820000 486.400000 ;
      RECT 281.620000 485.320000 324.820000 486.400000 ;
      RECT 236.620000 485.320000 279.820000 486.400000 ;
      RECT 191.620000 485.320000 234.820000 486.400000 ;
      RECT 146.620000 485.320000 189.820000 486.400000 ;
      RECT 101.620000 485.320000 144.820000 486.400000 ;
      RECT 56.620000 485.320000 99.820000 486.400000 ;
      RECT 11.620000 485.320000 54.820000 486.400000 ;
      RECT 4.860000 485.320000 9.655000 486.400000 ;
      RECT 0.000000 485.320000 3.060000 486.400000 ;
      RECT 0.000000 483.680000 550.160000 485.320000 ;
      RECT 544.900000 482.660000 550.160000 483.680000 ;
      RECT 544.900000 482.600000 548.960000 482.660000 ;
      RECT 508.620000 482.600000 543.100000 483.680000 ;
      RECT 463.620000 482.600000 506.820000 483.680000 ;
      RECT 418.620000 482.600000 461.820000 483.680000 ;
      RECT 373.620000 482.600000 416.820000 483.680000 ;
      RECT 328.620000 482.600000 371.820000 483.680000 ;
      RECT 283.620000 482.600000 326.820000 483.680000 ;
      RECT 238.620000 482.600000 281.820000 483.680000 ;
      RECT 193.620000 482.600000 236.820000 483.680000 ;
      RECT 148.620000 482.600000 191.820000 483.680000 ;
      RECT 103.620000 482.600000 146.820000 483.680000 ;
      RECT 58.620000 482.600000 101.820000 483.680000 ;
      RECT 13.620000 482.600000 56.820000 483.680000 ;
      RECT 7.060000 482.600000 11.820000 483.680000 ;
      RECT 0.000000 482.600000 5.260000 483.680000 ;
      RECT 0.000000 481.680000 548.960000 482.600000 ;
      RECT 0.000000 480.960000 550.160000 481.680000 ;
      RECT 547.100000 479.880000 550.160000 480.960000 ;
      RECT 506.620000 479.880000 545.300000 480.960000 ;
      RECT 461.620000 479.880000 504.820000 480.960000 ;
      RECT 416.620000 479.880000 459.820000 480.960000 ;
      RECT 371.620000 479.880000 414.820000 480.960000 ;
      RECT 326.620000 479.880000 369.820000 480.960000 ;
      RECT 281.620000 479.880000 324.820000 480.960000 ;
      RECT 236.620000 479.880000 279.820000 480.960000 ;
      RECT 191.620000 479.880000 234.820000 480.960000 ;
      RECT 146.620000 479.880000 189.820000 480.960000 ;
      RECT 101.620000 479.880000 144.820000 480.960000 ;
      RECT 56.620000 479.880000 99.820000 480.960000 ;
      RECT 11.620000 479.880000 54.820000 480.960000 ;
      RECT 4.860000 479.880000 9.655000 480.960000 ;
      RECT 0.000000 479.880000 3.060000 480.960000 ;
      RECT 0.000000 479.610000 550.160000 479.880000 ;
      RECT 0.000000 478.630000 548.960000 479.610000 ;
      RECT 0.000000 478.240000 550.160000 478.630000 ;
      RECT 544.900000 477.160000 550.160000 478.240000 ;
      RECT 508.620000 477.160000 543.100000 478.240000 ;
      RECT 463.620000 477.160000 506.820000 478.240000 ;
      RECT 418.620000 477.160000 461.820000 478.240000 ;
      RECT 373.620000 477.160000 416.820000 478.240000 ;
      RECT 328.620000 477.160000 371.820000 478.240000 ;
      RECT 283.620000 477.160000 326.820000 478.240000 ;
      RECT 238.620000 477.160000 281.820000 478.240000 ;
      RECT 193.620000 477.160000 236.820000 478.240000 ;
      RECT 148.620000 477.160000 191.820000 478.240000 ;
      RECT 103.620000 477.160000 146.820000 478.240000 ;
      RECT 58.620000 477.160000 101.820000 478.240000 ;
      RECT 13.620000 477.160000 56.820000 478.240000 ;
      RECT 7.060000 477.160000 11.820000 478.240000 ;
      RECT 0.000000 477.160000 5.260000 478.240000 ;
      RECT 0.000000 476.560000 550.160000 477.160000 ;
      RECT 0.000000 475.580000 548.960000 476.560000 ;
      RECT 0.000000 475.520000 550.160000 475.580000 ;
      RECT 547.100000 474.440000 550.160000 475.520000 ;
      RECT 506.620000 474.440000 545.300000 475.520000 ;
      RECT 461.620000 474.440000 504.820000 475.520000 ;
      RECT 416.620000 474.440000 459.820000 475.520000 ;
      RECT 371.620000 474.440000 414.820000 475.520000 ;
      RECT 326.620000 474.440000 369.820000 475.520000 ;
      RECT 281.620000 474.440000 324.820000 475.520000 ;
      RECT 236.620000 474.440000 279.820000 475.520000 ;
      RECT 191.620000 474.440000 234.820000 475.520000 ;
      RECT 146.620000 474.440000 189.820000 475.520000 ;
      RECT 101.620000 474.440000 144.820000 475.520000 ;
      RECT 56.620000 474.440000 99.820000 475.520000 ;
      RECT 11.620000 474.440000 54.820000 475.520000 ;
      RECT 4.860000 474.440000 9.655000 475.520000 ;
      RECT 0.000000 474.440000 3.060000 475.520000 ;
      RECT 0.000000 473.510000 550.160000 474.440000 ;
      RECT 0.000000 472.800000 548.960000 473.510000 ;
      RECT 544.900000 472.530000 548.960000 472.800000 ;
      RECT 544.900000 471.720000 550.160000 472.530000 ;
      RECT 508.620000 471.720000 543.100000 472.800000 ;
      RECT 463.620000 471.720000 506.820000 472.800000 ;
      RECT 418.620000 471.720000 461.820000 472.800000 ;
      RECT 373.620000 471.720000 416.820000 472.800000 ;
      RECT 328.620000 471.720000 371.820000 472.800000 ;
      RECT 283.620000 471.720000 326.820000 472.800000 ;
      RECT 238.620000 471.720000 281.820000 472.800000 ;
      RECT 193.620000 471.720000 236.820000 472.800000 ;
      RECT 148.620000 471.720000 191.820000 472.800000 ;
      RECT 103.620000 471.720000 146.820000 472.800000 ;
      RECT 58.620000 471.720000 101.820000 472.800000 ;
      RECT 13.620000 471.720000 56.820000 472.800000 ;
      RECT 7.060000 471.720000 11.820000 472.800000 ;
      RECT 0.000000 471.720000 5.260000 472.800000 ;
      RECT 0.000000 470.460000 550.160000 471.720000 ;
      RECT 0.000000 470.080000 548.960000 470.460000 ;
      RECT 547.100000 469.480000 548.960000 470.080000 ;
      RECT 547.100000 469.000000 550.160000 469.480000 ;
      RECT 506.620000 469.000000 545.300000 470.080000 ;
      RECT 461.620000 469.000000 504.820000 470.080000 ;
      RECT 416.620000 469.000000 459.820000 470.080000 ;
      RECT 371.620000 469.000000 414.820000 470.080000 ;
      RECT 326.620000 469.000000 369.820000 470.080000 ;
      RECT 281.620000 469.000000 324.820000 470.080000 ;
      RECT 236.620000 469.000000 279.820000 470.080000 ;
      RECT 191.620000 469.000000 234.820000 470.080000 ;
      RECT 146.620000 469.000000 189.820000 470.080000 ;
      RECT 101.620000 469.000000 144.820000 470.080000 ;
      RECT 56.620000 469.000000 99.820000 470.080000 ;
      RECT 11.620000 469.000000 54.820000 470.080000 ;
      RECT 4.860000 469.000000 9.655000 470.080000 ;
      RECT 0.000000 469.000000 3.060000 470.080000 ;
      RECT 0.000000 467.410000 550.160000 469.000000 ;
      RECT 0.000000 467.360000 548.960000 467.410000 ;
      RECT 544.900000 466.430000 548.960000 467.360000 ;
      RECT 544.900000 466.280000 550.160000 466.430000 ;
      RECT 508.620000 466.280000 543.100000 467.360000 ;
      RECT 463.620000 466.280000 506.820000 467.360000 ;
      RECT 418.620000 466.280000 461.820000 467.360000 ;
      RECT 373.620000 466.280000 416.820000 467.360000 ;
      RECT 328.620000 466.280000 371.820000 467.360000 ;
      RECT 283.620000 466.280000 326.820000 467.360000 ;
      RECT 238.620000 466.280000 281.820000 467.360000 ;
      RECT 193.620000 466.280000 236.820000 467.360000 ;
      RECT 148.620000 466.280000 191.820000 467.360000 ;
      RECT 103.620000 466.280000 146.820000 467.360000 ;
      RECT 58.620000 466.280000 101.820000 467.360000 ;
      RECT 13.620000 466.280000 56.820000 467.360000 ;
      RECT 7.060000 466.280000 11.820000 467.360000 ;
      RECT 0.000000 466.280000 5.260000 467.360000 ;
      RECT 0.000000 464.640000 550.160000 466.280000 ;
      RECT 547.100000 463.750000 550.160000 464.640000 ;
      RECT 547.100000 463.560000 548.960000 463.750000 ;
      RECT 506.620000 463.560000 545.300000 464.640000 ;
      RECT 461.620000 463.560000 504.820000 464.640000 ;
      RECT 416.620000 463.560000 459.820000 464.640000 ;
      RECT 371.620000 463.560000 414.820000 464.640000 ;
      RECT 326.620000 463.560000 369.820000 464.640000 ;
      RECT 281.620000 463.560000 324.820000 464.640000 ;
      RECT 236.620000 463.560000 279.820000 464.640000 ;
      RECT 191.620000 463.560000 234.820000 464.640000 ;
      RECT 146.620000 463.560000 189.820000 464.640000 ;
      RECT 101.620000 463.560000 144.820000 464.640000 ;
      RECT 56.620000 463.560000 99.820000 464.640000 ;
      RECT 11.620000 463.560000 54.820000 464.640000 ;
      RECT 4.860000 463.560000 9.655000 464.640000 ;
      RECT 0.000000 463.560000 3.060000 464.640000 ;
      RECT 0.000000 462.770000 548.960000 463.560000 ;
      RECT 0.000000 461.920000 550.160000 462.770000 ;
      RECT 544.900000 460.840000 550.160000 461.920000 ;
      RECT 508.620000 460.840000 543.100000 461.920000 ;
      RECT 463.620000 460.840000 506.820000 461.920000 ;
      RECT 418.620000 460.840000 461.820000 461.920000 ;
      RECT 373.620000 460.840000 416.820000 461.920000 ;
      RECT 328.620000 460.840000 371.820000 461.920000 ;
      RECT 283.620000 460.840000 326.820000 461.920000 ;
      RECT 238.620000 460.840000 281.820000 461.920000 ;
      RECT 193.620000 460.840000 236.820000 461.920000 ;
      RECT 148.620000 460.840000 191.820000 461.920000 ;
      RECT 103.620000 460.840000 146.820000 461.920000 ;
      RECT 58.620000 460.840000 101.820000 461.920000 ;
      RECT 13.620000 460.840000 56.820000 461.920000 ;
      RECT 7.060000 460.840000 11.820000 461.920000 ;
      RECT 0.000000 460.840000 5.260000 461.920000 ;
      RECT 0.000000 460.700000 550.160000 460.840000 ;
      RECT 0.000000 459.720000 548.960000 460.700000 ;
      RECT 0.000000 459.200000 550.160000 459.720000 ;
      RECT 547.100000 458.120000 550.160000 459.200000 ;
      RECT 506.620000 458.120000 545.300000 459.200000 ;
      RECT 461.620000 458.120000 504.820000 459.200000 ;
      RECT 416.620000 458.120000 459.820000 459.200000 ;
      RECT 371.620000 458.120000 414.820000 459.200000 ;
      RECT 326.620000 458.120000 369.820000 459.200000 ;
      RECT 281.620000 458.120000 324.820000 459.200000 ;
      RECT 236.620000 458.120000 279.820000 459.200000 ;
      RECT 191.620000 458.120000 234.820000 459.200000 ;
      RECT 146.620000 458.120000 189.820000 459.200000 ;
      RECT 101.620000 458.120000 144.820000 459.200000 ;
      RECT 56.620000 458.120000 99.820000 459.200000 ;
      RECT 11.620000 458.120000 54.820000 459.200000 ;
      RECT 4.860000 458.120000 9.655000 459.200000 ;
      RECT 0.000000 458.120000 3.060000 459.200000 ;
      RECT 0.000000 457.650000 550.160000 458.120000 ;
      RECT 0.000000 456.670000 548.960000 457.650000 ;
      RECT 0.000000 456.480000 550.160000 456.670000 ;
      RECT 544.900000 455.400000 550.160000 456.480000 ;
      RECT 508.620000 455.400000 543.100000 456.480000 ;
      RECT 463.620000 455.400000 506.820000 456.480000 ;
      RECT 418.620000 455.400000 461.820000 456.480000 ;
      RECT 373.620000 455.400000 416.820000 456.480000 ;
      RECT 328.620000 455.400000 371.820000 456.480000 ;
      RECT 283.620000 455.400000 326.820000 456.480000 ;
      RECT 238.620000 455.400000 281.820000 456.480000 ;
      RECT 193.620000 455.400000 236.820000 456.480000 ;
      RECT 148.620000 455.400000 191.820000 456.480000 ;
      RECT 103.620000 455.400000 146.820000 456.480000 ;
      RECT 58.620000 455.400000 101.820000 456.480000 ;
      RECT 13.620000 455.400000 56.820000 456.480000 ;
      RECT 7.060000 455.400000 11.820000 456.480000 ;
      RECT 0.000000 455.400000 5.260000 456.480000 ;
      RECT 0.000000 454.600000 550.160000 455.400000 ;
      RECT 0.000000 453.760000 548.960000 454.600000 ;
      RECT 547.100000 453.620000 548.960000 453.760000 ;
      RECT 547.100000 452.680000 550.160000 453.620000 ;
      RECT 506.620000 452.680000 545.300000 453.760000 ;
      RECT 461.620000 452.680000 504.820000 453.760000 ;
      RECT 416.620000 452.680000 459.820000 453.760000 ;
      RECT 371.620000 452.680000 414.820000 453.760000 ;
      RECT 326.620000 452.680000 369.820000 453.760000 ;
      RECT 281.620000 452.680000 324.820000 453.760000 ;
      RECT 236.620000 452.680000 279.820000 453.760000 ;
      RECT 191.620000 452.680000 234.820000 453.760000 ;
      RECT 146.620000 452.680000 189.820000 453.760000 ;
      RECT 101.620000 452.680000 144.820000 453.760000 ;
      RECT 56.620000 452.680000 99.820000 453.760000 ;
      RECT 11.620000 452.680000 54.820000 453.760000 ;
      RECT 4.860000 452.680000 9.655000 453.760000 ;
      RECT 0.000000 452.680000 3.060000 453.760000 ;
      RECT 0.000000 451.550000 550.160000 452.680000 ;
      RECT 0.000000 451.040000 548.960000 451.550000 ;
      RECT 544.900000 450.570000 548.960000 451.040000 ;
      RECT 544.900000 449.960000 550.160000 450.570000 ;
      RECT 508.620000 449.960000 543.100000 451.040000 ;
      RECT 463.620000 449.960000 506.820000 451.040000 ;
      RECT 418.620000 449.960000 461.820000 451.040000 ;
      RECT 373.620000 449.960000 416.820000 451.040000 ;
      RECT 328.620000 449.960000 371.820000 451.040000 ;
      RECT 283.620000 449.960000 326.820000 451.040000 ;
      RECT 238.620000 449.960000 281.820000 451.040000 ;
      RECT 193.620000 449.960000 236.820000 451.040000 ;
      RECT 148.620000 449.960000 191.820000 451.040000 ;
      RECT 103.620000 449.960000 146.820000 451.040000 ;
      RECT 58.620000 449.960000 101.820000 451.040000 ;
      RECT 13.620000 449.960000 56.820000 451.040000 ;
      RECT 7.060000 449.960000 11.820000 451.040000 ;
      RECT 0.000000 449.960000 5.260000 451.040000 ;
      RECT 0.000000 448.500000 550.160000 449.960000 ;
      RECT 0.000000 448.320000 548.960000 448.500000 ;
      RECT 547.100000 447.520000 548.960000 448.320000 ;
      RECT 547.100000 447.240000 550.160000 447.520000 ;
      RECT 506.620000 447.240000 545.300000 448.320000 ;
      RECT 461.620000 447.240000 504.820000 448.320000 ;
      RECT 416.620000 447.240000 459.820000 448.320000 ;
      RECT 371.620000 447.240000 414.820000 448.320000 ;
      RECT 326.620000 447.240000 369.820000 448.320000 ;
      RECT 281.620000 447.240000 324.820000 448.320000 ;
      RECT 236.620000 447.240000 279.820000 448.320000 ;
      RECT 191.620000 447.240000 234.820000 448.320000 ;
      RECT 146.620000 447.240000 189.820000 448.320000 ;
      RECT 101.620000 447.240000 144.820000 448.320000 ;
      RECT 56.620000 447.240000 99.820000 448.320000 ;
      RECT 11.620000 447.240000 54.820000 448.320000 ;
      RECT 4.860000 447.240000 9.655000 448.320000 ;
      RECT 0.000000 447.240000 3.060000 448.320000 ;
      RECT 0.000000 445.600000 550.160000 447.240000 ;
      RECT 544.900000 444.840000 550.160000 445.600000 ;
      RECT 544.900000 444.520000 548.960000 444.840000 ;
      RECT 508.620000 444.520000 543.100000 445.600000 ;
      RECT 463.620000 444.520000 506.820000 445.600000 ;
      RECT 418.620000 444.520000 461.820000 445.600000 ;
      RECT 373.620000 444.520000 416.820000 445.600000 ;
      RECT 328.620000 444.520000 371.820000 445.600000 ;
      RECT 283.620000 444.520000 326.820000 445.600000 ;
      RECT 238.620000 444.520000 281.820000 445.600000 ;
      RECT 193.620000 444.520000 236.820000 445.600000 ;
      RECT 148.620000 444.520000 191.820000 445.600000 ;
      RECT 103.620000 444.520000 146.820000 445.600000 ;
      RECT 58.620000 444.520000 101.820000 445.600000 ;
      RECT 13.620000 444.520000 56.820000 445.600000 ;
      RECT 7.060000 444.520000 11.820000 445.600000 ;
      RECT 0.000000 444.520000 5.260000 445.600000 ;
      RECT 0.000000 443.860000 548.960000 444.520000 ;
      RECT 0.000000 442.880000 550.160000 443.860000 ;
      RECT 547.100000 441.800000 550.160000 442.880000 ;
      RECT 506.620000 441.800000 545.300000 442.880000 ;
      RECT 461.620000 441.800000 504.820000 442.880000 ;
      RECT 416.620000 441.800000 459.820000 442.880000 ;
      RECT 371.620000 441.800000 414.820000 442.880000 ;
      RECT 326.620000 441.800000 369.820000 442.880000 ;
      RECT 281.620000 441.800000 324.820000 442.880000 ;
      RECT 236.620000 441.800000 279.820000 442.880000 ;
      RECT 191.620000 441.800000 234.820000 442.880000 ;
      RECT 146.620000 441.800000 189.820000 442.880000 ;
      RECT 101.620000 441.800000 144.820000 442.880000 ;
      RECT 56.620000 441.800000 99.820000 442.880000 ;
      RECT 11.620000 441.800000 54.820000 442.880000 ;
      RECT 4.860000 441.800000 9.655000 442.880000 ;
      RECT 0.000000 441.800000 3.060000 442.880000 ;
      RECT 0.000000 441.790000 550.160000 441.800000 ;
      RECT 0.000000 440.810000 548.960000 441.790000 ;
      RECT 0.000000 440.160000 550.160000 440.810000 ;
      RECT 544.900000 439.080000 550.160000 440.160000 ;
      RECT 508.620000 439.080000 543.100000 440.160000 ;
      RECT 463.620000 439.080000 506.820000 440.160000 ;
      RECT 418.620000 439.080000 461.820000 440.160000 ;
      RECT 373.620000 439.080000 416.820000 440.160000 ;
      RECT 328.620000 439.080000 371.820000 440.160000 ;
      RECT 283.620000 439.080000 326.820000 440.160000 ;
      RECT 238.620000 439.080000 281.820000 440.160000 ;
      RECT 193.620000 439.080000 236.820000 440.160000 ;
      RECT 148.620000 439.080000 191.820000 440.160000 ;
      RECT 103.620000 439.080000 146.820000 440.160000 ;
      RECT 58.620000 439.080000 101.820000 440.160000 ;
      RECT 13.620000 439.080000 56.820000 440.160000 ;
      RECT 7.060000 439.080000 11.820000 440.160000 ;
      RECT 0.000000 439.080000 5.260000 440.160000 ;
      RECT 0.000000 438.740000 550.160000 439.080000 ;
      RECT 0.000000 437.760000 548.960000 438.740000 ;
      RECT 0.000000 437.440000 550.160000 437.760000 ;
      RECT 547.100000 436.360000 550.160000 437.440000 ;
      RECT 506.620000 436.360000 545.300000 437.440000 ;
      RECT 461.620000 436.360000 504.820000 437.440000 ;
      RECT 416.620000 436.360000 459.820000 437.440000 ;
      RECT 371.620000 436.360000 414.820000 437.440000 ;
      RECT 326.620000 436.360000 369.820000 437.440000 ;
      RECT 281.620000 436.360000 324.820000 437.440000 ;
      RECT 236.620000 436.360000 279.820000 437.440000 ;
      RECT 191.620000 436.360000 234.820000 437.440000 ;
      RECT 146.620000 436.360000 189.820000 437.440000 ;
      RECT 101.620000 436.360000 144.820000 437.440000 ;
      RECT 56.620000 436.360000 99.820000 437.440000 ;
      RECT 11.620000 436.360000 54.820000 437.440000 ;
      RECT 4.860000 436.360000 9.655000 437.440000 ;
      RECT 0.000000 436.360000 3.060000 437.440000 ;
      RECT 0.000000 435.690000 550.160000 436.360000 ;
      RECT 0.000000 434.720000 548.960000 435.690000 ;
      RECT 544.900000 434.710000 548.960000 434.720000 ;
      RECT 544.900000 433.640000 550.160000 434.710000 ;
      RECT 508.620000 433.640000 543.100000 434.720000 ;
      RECT 463.620000 433.640000 506.820000 434.720000 ;
      RECT 418.620000 433.640000 461.820000 434.720000 ;
      RECT 373.620000 433.640000 416.820000 434.720000 ;
      RECT 328.620000 433.640000 371.820000 434.720000 ;
      RECT 283.620000 433.640000 326.820000 434.720000 ;
      RECT 238.620000 433.640000 281.820000 434.720000 ;
      RECT 193.620000 433.640000 236.820000 434.720000 ;
      RECT 148.620000 433.640000 191.820000 434.720000 ;
      RECT 103.620000 433.640000 146.820000 434.720000 ;
      RECT 58.620000 433.640000 101.820000 434.720000 ;
      RECT 13.620000 433.640000 56.820000 434.720000 ;
      RECT 7.060000 433.640000 11.820000 434.720000 ;
      RECT 0.000000 433.640000 5.260000 434.720000 ;
      RECT 0.000000 432.640000 550.160000 433.640000 ;
      RECT 0.000000 432.000000 548.960000 432.640000 ;
      RECT 547.100000 431.660000 548.960000 432.000000 ;
      RECT 547.100000 430.920000 550.160000 431.660000 ;
      RECT 506.620000 430.920000 545.300000 432.000000 ;
      RECT 461.620000 430.920000 504.820000 432.000000 ;
      RECT 416.620000 430.920000 459.820000 432.000000 ;
      RECT 371.620000 430.920000 414.820000 432.000000 ;
      RECT 326.620000 430.920000 369.820000 432.000000 ;
      RECT 281.620000 430.920000 324.820000 432.000000 ;
      RECT 236.620000 430.920000 279.820000 432.000000 ;
      RECT 191.620000 430.920000 234.820000 432.000000 ;
      RECT 146.620000 430.920000 189.820000 432.000000 ;
      RECT 101.620000 430.920000 144.820000 432.000000 ;
      RECT 56.620000 430.920000 99.820000 432.000000 ;
      RECT 11.620000 430.920000 54.820000 432.000000 ;
      RECT 4.860000 430.920000 9.655000 432.000000 ;
      RECT 0.000000 430.920000 3.060000 432.000000 ;
      RECT 0.000000 429.590000 550.160000 430.920000 ;
      RECT 0.000000 429.280000 548.960000 429.590000 ;
      RECT 544.900000 428.610000 548.960000 429.280000 ;
      RECT 544.900000 428.200000 550.160000 428.610000 ;
      RECT 508.620000 428.200000 543.100000 429.280000 ;
      RECT 463.620000 428.200000 506.820000 429.280000 ;
      RECT 418.620000 428.200000 461.820000 429.280000 ;
      RECT 373.620000 428.200000 416.820000 429.280000 ;
      RECT 328.620000 428.200000 371.820000 429.280000 ;
      RECT 283.620000 428.200000 326.820000 429.280000 ;
      RECT 238.620000 428.200000 281.820000 429.280000 ;
      RECT 193.620000 428.200000 236.820000 429.280000 ;
      RECT 148.620000 428.200000 191.820000 429.280000 ;
      RECT 103.620000 428.200000 146.820000 429.280000 ;
      RECT 58.620000 428.200000 101.820000 429.280000 ;
      RECT 13.620000 428.200000 56.820000 429.280000 ;
      RECT 7.060000 428.200000 11.820000 429.280000 ;
      RECT 0.000000 428.200000 5.260000 429.280000 ;
      RECT 0.000000 426.560000 550.160000 428.200000 ;
      RECT 547.100000 425.930000 550.160000 426.560000 ;
      RECT 547.100000 425.480000 548.960000 425.930000 ;
      RECT 506.620000 425.480000 545.300000 426.560000 ;
      RECT 461.620000 425.480000 504.820000 426.560000 ;
      RECT 416.620000 425.480000 459.820000 426.560000 ;
      RECT 371.620000 425.480000 414.820000 426.560000 ;
      RECT 326.620000 425.480000 369.820000 426.560000 ;
      RECT 281.620000 425.480000 324.820000 426.560000 ;
      RECT 236.620000 425.480000 279.820000 426.560000 ;
      RECT 191.620000 425.480000 234.820000 426.560000 ;
      RECT 146.620000 425.480000 189.820000 426.560000 ;
      RECT 101.620000 425.480000 144.820000 426.560000 ;
      RECT 56.620000 425.480000 99.820000 426.560000 ;
      RECT 11.620000 425.480000 54.820000 426.560000 ;
      RECT 4.860000 425.480000 9.655000 426.560000 ;
      RECT 0.000000 425.480000 3.060000 426.560000 ;
      RECT 0.000000 424.950000 548.960000 425.480000 ;
      RECT 0.000000 423.840000 550.160000 424.950000 ;
      RECT 544.900000 422.880000 550.160000 423.840000 ;
      RECT 544.900000 422.760000 548.960000 422.880000 ;
      RECT 508.620000 422.760000 543.100000 423.840000 ;
      RECT 463.620000 422.760000 506.820000 423.840000 ;
      RECT 418.620000 422.760000 461.820000 423.840000 ;
      RECT 373.620000 422.760000 416.820000 423.840000 ;
      RECT 328.620000 422.760000 371.820000 423.840000 ;
      RECT 283.620000 422.760000 326.820000 423.840000 ;
      RECT 238.620000 422.760000 281.820000 423.840000 ;
      RECT 193.620000 422.760000 236.820000 423.840000 ;
      RECT 148.620000 422.760000 191.820000 423.840000 ;
      RECT 103.620000 422.760000 146.820000 423.840000 ;
      RECT 58.620000 422.760000 101.820000 423.840000 ;
      RECT 13.620000 422.760000 56.820000 423.840000 ;
      RECT 7.060000 422.760000 11.820000 423.840000 ;
      RECT 0.000000 422.760000 5.260000 423.840000 ;
      RECT 0.000000 421.900000 548.960000 422.760000 ;
      RECT 0.000000 421.120000 550.160000 421.900000 ;
      RECT 547.100000 420.040000 550.160000 421.120000 ;
      RECT 506.620000 420.040000 545.300000 421.120000 ;
      RECT 461.620000 420.040000 504.820000 421.120000 ;
      RECT 416.620000 420.040000 459.820000 421.120000 ;
      RECT 371.620000 420.040000 414.820000 421.120000 ;
      RECT 326.620000 420.040000 369.820000 421.120000 ;
      RECT 281.620000 420.040000 324.820000 421.120000 ;
      RECT 236.620000 420.040000 279.820000 421.120000 ;
      RECT 191.620000 420.040000 234.820000 421.120000 ;
      RECT 146.620000 420.040000 189.820000 421.120000 ;
      RECT 101.620000 420.040000 144.820000 421.120000 ;
      RECT 56.620000 420.040000 99.820000 421.120000 ;
      RECT 11.620000 420.040000 54.820000 421.120000 ;
      RECT 4.860000 420.040000 9.655000 421.120000 ;
      RECT 0.000000 420.040000 3.060000 421.120000 ;
      RECT 0.000000 419.830000 550.160000 420.040000 ;
      RECT 0.000000 418.850000 548.960000 419.830000 ;
      RECT 0.000000 418.400000 550.160000 418.850000 ;
      RECT 544.900000 417.320000 550.160000 418.400000 ;
      RECT 508.620000 417.320000 543.100000 418.400000 ;
      RECT 463.620000 417.320000 506.820000 418.400000 ;
      RECT 418.620000 417.320000 461.820000 418.400000 ;
      RECT 373.620000 417.320000 416.820000 418.400000 ;
      RECT 328.620000 417.320000 371.820000 418.400000 ;
      RECT 283.620000 417.320000 326.820000 418.400000 ;
      RECT 238.620000 417.320000 281.820000 418.400000 ;
      RECT 193.620000 417.320000 236.820000 418.400000 ;
      RECT 148.620000 417.320000 191.820000 418.400000 ;
      RECT 103.620000 417.320000 146.820000 418.400000 ;
      RECT 58.620000 417.320000 101.820000 418.400000 ;
      RECT 13.620000 417.320000 56.820000 418.400000 ;
      RECT 7.060000 417.320000 11.820000 418.400000 ;
      RECT 0.000000 417.320000 5.260000 418.400000 ;
      RECT 0.000000 416.780000 550.160000 417.320000 ;
      RECT 0.000000 415.800000 548.960000 416.780000 ;
      RECT 0.000000 415.680000 550.160000 415.800000 ;
      RECT 547.100000 414.600000 550.160000 415.680000 ;
      RECT 506.620000 414.600000 545.300000 415.680000 ;
      RECT 461.620000 414.600000 504.820000 415.680000 ;
      RECT 416.620000 414.600000 459.820000 415.680000 ;
      RECT 371.620000 414.600000 414.820000 415.680000 ;
      RECT 326.620000 414.600000 369.820000 415.680000 ;
      RECT 281.620000 414.600000 324.820000 415.680000 ;
      RECT 236.620000 414.600000 279.820000 415.680000 ;
      RECT 191.620000 414.600000 234.820000 415.680000 ;
      RECT 146.620000 414.600000 189.820000 415.680000 ;
      RECT 101.620000 414.600000 144.820000 415.680000 ;
      RECT 56.620000 414.600000 99.820000 415.680000 ;
      RECT 11.620000 414.600000 54.820000 415.680000 ;
      RECT 4.860000 414.600000 9.655000 415.680000 ;
      RECT 0.000000 414.600000 3.060000 415.680000 ;
      RECT 0.000000 413.730000 550.160000 414.600000 ;
      RECT 0.000000 412.960000 548.960000 413.730000 ;
      RECT 544.900000 412.750000 548.960000 412.960000 ;
      RECT 544.900000 411.880000 550.160000 412.750000 ;
      RECT 508.620000 411.880000 543.100000 412.960000 ;
      RECT 463.620000 411.880000 506.820000 412.960000 ;
      RECT 418.620000 411.880000 461.820000 412.960000 ;
      RECT 373.620000 411.880000 416.820000 412.960000 ;
      RECT 328.620000 411.880000 371.820000 412.960000 ;
      RECT 283.620000 411.880000 326.820000 412.960000 ;
      RECT 238.620000 411.880000 281.820000 412.960000 ;
      RECT 193.620000 411.880000 236.820000 412.960000 ;
      RECT 148.620000 411.880000 191.820000 412.960000 ;
      RECT 103.620000 411.880000 146.820000 412.960000 ;
      RECT 58.620000 411.880000 101.820000 412.960000 ;
      RECT 13.620000 411.880000 56.820000 412.960000 ;
      RECT 7.060000 411.880000 11.820000 412.960000 ;
      RECT 0.000000 411.880000 5.260000 412.960000 ;
      RECT 0.000000 410.680000 550.160000 411.880000 ;
      RECT 0.000000 410.240000 548.960000 410.680000 ;
      RECT 547.100000 409.700000 548.960000 410.240000 ;
      RECT 547.100000 409.160000 550.160000 409.700000 ;
      RECT 506.620000 409.160000 545.300000 410.240000 ;
      RECT 461.620000 409.160000 504.820000 410.240000 ;
      RECT 416.620000 409.160000 459.820000 410.240000 ;
      RECT 371.620000 409.160000 414.820000 410.240000 ;
      RECT 326.620000 409.160000 369.820000 410.240000 ;
      RECT 281.620000 409.160000 324.820000 410.240000 ;
      RECT 236.620000 409.160000 279.820000 410.240000 ;
      RECT 191.620000 409.160000 234.820000 410.240000 ;
      RECT 146.620000 409.160000 189.820000 410.240000 ;
      RECT 101.620000 409.160000 144.820000 410.240000 ;
      RECT 56.620000 409.160000 99.820000 410.240000 ;
      RECT 11.620000 409.160000 54.820000 410.240000 ;
      RECT 4.860000 409.160000 9.655000 410.240000 ;
      RECT 0.000000 409.160000 3.060000 410.240000 ;
      RECT 0.000000 407.520000 550.160000 409.160000 ;
      RECT 544.900000 407.020000 550.160000 407.520000 ;
      RECT 544.900000 406.440000 548.960000 407.020000 ;
      RECT 508.620000 406.440000 543.100000 407.520000 ;
      RECT 463.620000 406.440000 506.820000 407.520000 ;
      RECT 418.620000 406.440000 461.820000 407.520000 ;
      RECT 373.620000 406.440000 416.820000 407.520000 ;
      RECT 328.620000 406.440000 371.820000 407.520000 ;
      RECT 283.620000 406.440000 326.820000 407.520000 ;
      RECT 238.620000 406.440000 281.820000 407.520000 ;
      RECT 193.620000 406.440000 236.820000 407.520000 ;
      RECT 148.620000 406.440000 191.820000 407.520000 ;
      RECT 103.620000 406.440000 146.820000 407.520000 ;
      RECT 58.620000 406.440000 101.820000 407.520000 ;
      RECT 13.620000 406.440000 56.820000 407.520000 ;
      RECT 7.060000 406.440000 11.820000 407.520000 ;
      RECT 0.000000 406.440000 5.260000 407.520000 ;
      RECT 0.000000 406.040000 548.960000 406.440000 ;
      RECT 0.000000 404.800000 550.160000 406.040000 ;
      RECT 547.100000 403.970000 550.160000 404.800000 ;
      RECT 547.100000 403.720000 548.960000 403.970000 ;
      RECT 506.620000 403.720000 545.300000 404.800000 ;
      RECT 461.620000 403.720000 504.820000 404.800000 ;
      RECT 416.620000 403.720000 459.820000 404.800000 ;
      RECT 371.620000 403.720000 414.820000 404.800000 ;
      RECT 326.620000 403.720000 369.820000 404.800000 ;
      RECT 281.620000 403.720000 324.820000 404.800000 ;
      RECT 236.620000 403.720000 279.820000 404.800000 ;
      RECT 191.620000 403.720000 234.820000 404.800000 ;
      RECT 146.620000 403.720000 189.820000 404.800000 ;
      RECT 101.620000 403.720000 144.820000 404.800000 ;
      RECT 56.620000 403.720000 99.820000 404.800000 ;
      RECT 11.620000 403.720000 54.820000 404.800000 ;
      RECT 4.860000 403.720000 9.655000 404.800000 ;
      RECT 0.000000 403.720000 3.060000 404.800000 ;
      RECT 0.000000 402.990000 548.960000 403.720000 ;
      RECT 0.000000 402.080000 550.160000 402.990000 ;
      RECT 544.900000 401.000000 550.160000 402.080000 ;
      RECT 508.620000 401.000000 543.100000 402.080000 ;
      RECT 463.620000 401.000000 506.820000 402.080000 ;
      RECT 418.620000 401.000000 461.820000 402.080000 ;
      RECT 373.620000 401.000000 416.820000 402.080000 ;
      RECT 328.620000 401.000000 371.820000 402.080000 ;
      RECT 283.620000 401.000000 326.820000 402.080000 ;
      RECT 238.620000 401.000000 281.820000 402.080000 ;
      RECT 193.620000 401.000000 236.820000 402.080000 ;
      RECT 148.620000 401.000000 191.820000 402.080000 ;
      RECT 103.620000 401.000000 146.820000 402.080000 ;
      RECT 58.620000 401.000000 101.820000 402.080000 ;
      RECT 13.620000 401.000000 56.820000 402.080000 ;
      RECT 7.060000 401.000000 11.820000 402.080000 ;
      RECT 0.000000 401.000000 5.260000 402.080000 ;
      RECT 0.000000 400.920000 550.160000 401.000000 ;
      RECT 0.000000 399.940000 548.960000 400.920000 ;
      RECT 0.000000 399.360000 550.160000 399.940000 ;
      RECT 547.100000 398.280000 550.160000 399.360000 ;
      RECT 506.620000 398.280000 545.300000 399.360000 ;
      RECT 461.620000 398.280000 504.820000 399.360000 ;
      RECT 416.620000 398.280000 459.820000 399.360000 ;
      RECT 371.620000 398.280000 414.820000 399.360000 ;
      RECT 326.620000 398.280000 369.820000 399.360000 ;
      RECT 281.620000 398.280000 324.820000 399.360000 ;
      RECT 236.620000 398.280000 279.820000 399.360000 ;
      RECT 191.620000 398.280000 234.820000 399.360000 ;
      RECT 146.620000 398.280000 189.820000 399.360000 ;
      RECT 101.620000 398.280000 144.820000 399.360000 ;
      RECT 56.620000 398.280000 99.820000 399.360000 ;
      RECT 11.620000 398.280000 54.820000 399.360000 ;
      RECT 4.860000 398.280000 9.655000 399.360000 ;
      RECT 0.000000 398.280000 3.060000 399.360000 ;
      RECT 0.000000 397.870000 550.160000 398.280000 ;
      RECT 0.000000 396.890000 548.960000 397.870000 ;
      RECT 0.000000 396.640000 550.160000 396.890000 ;
      RECT 544.900000 395.560000 550.160000 396.640000 ;
      RECT 508.620000 395.560000 543.100000 396.640000 ;
      RECT 463.620000 395.560000 506.820000 396.640000 ;
      RECT 418.620000 395.560000 461.820000 396.640000 ;
      RECT 373.620000 395.560000 416.820000 396.640000 ;
      RECT 328.620000 395.560000 371.820000 396.640000 ;
      RECT 283.620000 395.560000 326.820000 396.640000 ;
      RECT 238.620000 395.560000 281.820000 396.640000 ;
      RECT 193.620000 395.560000 236.820000 396.640000 ;
      RECT 148.620000 395.560000 191.820000 396.640000 ;
      RECT 103.620000 395.560000 146.820000 396.640000 ;
      RECT 58.620000 395.560000 101.820000 396.640000 ;
      RECT 13.620000 395.560000 56.820000 396.640000 ;
      RECT 7.060000 395.560000 11.820000 396.640000 ;
      RECT 0.000000 395.560000 5.260000 396.640000 ;
      RECT 0.000000 394.820000 550.160000 395.560000 ;
      RECT 0.000000 393.920000 548.960000 394.820000 ;
      RECT 547.100000 393.840000 548.960000 393.920000 ;
      RECT 547.100000 392.840000 550.160000 393.840000 ;
      RECT 506.620000 392.840000 545.300000 393.920000 ;
      RECT 461.620000 392.840000 504.820000 393.920000 ;
      RECT 416.620000 392.840000 459.820000 393.920000 ;
      RECT 371.620000 392.840000 414.820000 393.920000 ;
      RECT 326.620000 392.840000 369.820000 393.920000 ;
      RECT 281.620000 392.840000 324.820000 393.920000 ;
      RECT 236.620000 392.840000 279.820000 393.920000 ;
      RECT 191.620000 392.840000 234.820000 393.920000 ;
      RECT 146.620000 392.840000 189.820000 393.920000 ;
      RECT 101.620000 392.840000 144.820000 393.920000 ;
      RECT 56.620000 392.840000 99.820000 393.920000 ;
      RECT 11.620000 392.840000 54.820000 393.920000 ;
      RECT 4.860000 392.840000 9.655000 393.920000 ;
      RECT 0.000000 392.840000 3.060000 393.920000 ;
      RECT 0.000000 391.770000 550.160000 392.840000 ;
      RECT 0.000000 391.200000 548.960000 391.770000 ;
      RECT 544.900000 390.790000 548.960000 391.200000 ;
      RECT 544.900000 390.120000 550.160000 390.790000 ;
      RECT 508.620000 390.120000 543.100000 391.200000 ;
      RECT 463.620000 390.120000 506.820000 391.200000 ;
      RECT 418.620000 390.120000 461.820000 391.200000 ;
      RECT 373.620000 390.120000 416.820000 391.200000 ;
      RECT 328.620000 390.120000 371.820000 391.200000 ;
      RECT 283.620000 390.120000 326.820000 391.200000 ;
      RECT 238.620000 390.120000 281.820000 391.200000 ;
      RECT 193.620000 390.120000 236.820000 391.200000 ;
      RECT 148.620000 390.120000 191.820000 391.200000 ;
      RECT 103.620000 390.120000 146.820000 391.200000 ;
      RECT 58.620000 390.120000 101.820000 391.200000 ;
      RECT 13.620000 390.120000 56.820000 391.200000 ;
      RECT 7.060000 390.120000 11.820000 391.200000 ;
      RECT 0.000000 390.120000 5.260000 391.200000 ;
      RECT 0.000000 388.720000 550.160000 390.120000 ;
      RECT 0.000000 388.480000 548.960000 388.720000 ;
      RECT 547.100000 387.740000 548.960000 388.480000 ;
      RECT 547.100000 387.400000 550.160000 387.740000 ;
      RECT 506.620000 387.400000 545.300000 388.480000 ;
      RECT 461.620000 387.400000 504.820000 388.480000 ;
      RECT 416.620000 387.400000 459.820000 388.480000 ;
      RECT 371.620000 387.400000 414.820000 388.480000 ;
      RECT 326.620000 387.400000 369.820000 388.480000 ;
      RECT 281.620000 387.400000 324.820000 388.480000 ;
      RECT 236.620000 387.400000 279.820000 388.480000 ;
      RECT 191.620000 387.400000 234.820000 388.480000 ;
      RECT 146.620000 387.400000 189.820000 388.480000 ;
      RECT 101.620000 387.400000 144.820000 388.480000 ;
      RECT 56.620000 387.400000 99.820000 388.480000 ;
      RECT 11.620000 387.400000 54.820000 388.480000 ;
      RECT 4.860000 387.400000 9.655000 388.480000 ;
      RECT 0.000000 387.400000 3.060000 388.480000 ;
      RECT 0.000000 385.760000 550.160000 387.400000 ;
      RECT 544.900000 385.060000 550.160000 385.760000 ;
      RECT 544.900000 384.680000 548.960000 385.060000 ;
      RECT 508.620000 384.680000 543.100000 385.760000 ;
      RECT 463.620000 384.680000 506.820000 385.760000 ;
      RECT 418.620000 384.680000 461.820000 385.760000 ;
      RECT 373.620000 384.680000 416.820000 385.760000 ;
      RECT 328.620000 384.680000 371.820000 385.760000 ;
      RECT 283.620000 384.680000 326.820000 385.760000 ;
      RECT 238.620000 384.680000 281.820000 385.760000 ;
      RECT 193.620000 384.680000 236.820000 385.760000 ;
      RECT 148.620000 384.680000 191.820000 385.760000 ;
      RECT 103.620000 384.680000 146.820000 385.760000 ;
      RECT 58.620000 384.680000 101.820000 385.760000 ;
      RECT 13.620000 384.680000 56.820000 385.760000 ;
      RECT 7.060000 384.680000 11.820000 385.760000 ;
      RECT 0.000000 384.680000 5.260000 385.760000 ;
      RECT 0.000000 384.080000 548.960000 384.680000 ;
      RECT 0.000000 383.040000 550.160000 384.080000 ;
      RECT 547.100000 382.010000 550.160000 383.040000 ;
      RECT 547.100000 381.960000 548.960000 382.010000 ;
      RECT 506.620000 381.960000 545.300000 383.040000 ;
      RECT 461.620000 381.960000 504.820000 383.040000 ;
      RECT 416.620000 381.960000 459.820000 383.040000 ;
      RECT 371.620000 381.960000 414.820000 383.040000 ;
      RECT 326.620000 381.960000 369.820000 383.040000 ;
      RECT 281.620000 381.960000 324.820000 383.040000 ;
      RECT 236.620000 381.960000 279.820000 383.040000 ;
      RECT 191.620000 381.960000 234.820000 383.040000 ;
      RECT 146.620000 381.960000 189.820000 383.040000 ;
      RECT 101.620000 381.960000 144.820000 383.040000 ;
      RECT 56.620000 381.960000 99.820000 383.040000 ;
      RECT 11.620000 381.960000 54.820000 383.040000 ;
      RECT 4.860000 381.960000 9.655000 383.040000 ;
      RECT 0.000000 381.960000 3.060000 383.040000 ;
      RECT 0.000000 381.030000 548.960000 381.960000 ;
      RECT 0.000000 380.320000 550.160000 381.030000 ;
      RECT 544.900000 379.240000 550.160000 380.320000 ;
      RECT 508.620000 379.240000 543.100000 380.320000 ;
      RECT 463.620000 379.240000 506.820000 380.320000 ;
      RECT 418.620000 379.240000 461.820000 380.320000 ;
      RECT 373.620000 379.240000 416.820000 380.320000 ;
      RECT 328.620000 379.240000 371.820000 380.320000 ;
      RECT 283.620000 379.240000 326.820000 380.320000 ;
      RECT 238.620000 379.240000 281.820000 380.320000 ;
      RECT 193.620000 379.240000 236.820000 380.320000 ;
      RECT 148.620000 379.240000 191.820000 380.320000 ;
      RECT 103.620000 379.240000 146.820000 380.320000 ;
      RECT 58.620000 379.240000 101.820000 380.320000 ;
      RECT 13.620000 379.240000 56.820000 380.320000 ;
      RECT 7.060000 379.240000 11.820000 380.320000 ;
      RECT 0.000000 379.240000 5.260000 380.320000 ;
      RECT 0.000000 378.960000 550.160000 379.240000 ;
      RECT 0.000000 377.980000 548.960000 378.960000 ;
      RECT 0.000000 377.600000 550.160000 377.980000 ;
      RECT 547.100000 376.520000 550.160000 377.600000 ;
      RECT 506.620000 376.520000 545.300000 377.600000 ;
      RECT 461.620000 376.520000 504.820000 377.600000 ;
      RECT 416.620000 376.520000 459.820000 377.600000 ;
      RECT 371.620000 376.520000 414.820000 377.600000 ;
      RECT 326.620000 376.520000 369.820000 377.600000 ;
      RECT 281.620000 376.520000 324.820000 377.600000 ;
      RECT 236.620000 376.520000 279.820000 377.600000 ;
      RECT 191.620000 376.520000 234.820000 377.600000 ;
      RECT 146.620000 376.520000 189.820000 377.600000 ;
      RECT 101.620000 376.520000 144.820000 377.600000 ;
      RECT 56.620000 376.520000 99.820000 377.600000 ;
      RECT 11.620000 376.520000 54.820000 377.600000 ;
      RECT 4.860000 376.520000 9.655000 377.600000 ;
      RECT 0.000000 376.520000 3.060000 377.600000 ;
      RECT 0.000000 375.910000 550.160000 376.520000 ;
      RECT 0.000000 374.930000 548.960000 375.910000 ;
      RECT 0.000000 374.880000 550.160000 374.930000 ;
      RECT 544.900000 373.800000 550.160000 374.880000 ;
      RECT 508.620000 373.800000 543.100000 374.880000 ;
      RECT 463.620000 373.800000 506.820000 374.880000 ;
      RECT 418.620000 373.800000 461.820000 374.880000 ;
      RECT 373.620000 373.800000 416.820000 374.880000 ;
      RECT 328.620000 373.800000 371.820000 374.880000 ;
      RECT 283.620000 373.800000 326.820000 374.880000 ;
      RECT 238.620000 373.800000 281.820000 374.880000 ;
      RECT 193.620000 373.800000 236.820000 374.880000 ;
      RECT 148.620000 373.800000 191.820000 374.880000 ;
      RECT 103.620000 373.800000 146.820000 374.880000 ;
      RECT 58.620000 373.800000 101.820000 374.880000 ;
      RECT 13.620000 373.800000 56.820000 374.880000 ;
      RECT 7.060000 373.800000 11.820000 374.880000 ;
      RECT 0.000000 373.800000 5.260000 374.880000 ;
      RECT 0.000000 372.860000 550.160000 373.800000 ;
      RECT 0.000000 372.160000 548.960000 372.860000 ;
      RECT 547.100000 371.880000 548.960000 372.160000 ;
      RECT 547.100000 371.080000 550.160000 371.880000 ;
      RECT 506.620000 371.080000 545.300000 372.160000 ;
      RECT 461.620000 371.080000 504.820000 372.160000 ;
      RECT 416.620000 371.080000 459.820000 372.160000 ;
      RECT 371.620000 371.080000 414.820000 372.160000 ;
      RECT 326.620000 371.080000 369.820000 372.160000 ;
      RECT 281.620000 371.080000 324.820000 372.160000 ;
      RECT 236.620000 371.080000 279.820000 372.160000 ;
      RECT 191.620000 371.080000 234.820000 372.160000 ;
      RECT 146.620000 371.080000 189.820000 372.160000 ;
      RECT 101.620000 371.080000 144.820000 372.160000 ;
      RECT 56.620000 371.080000 99.820000 372.160000 ;
      RECT 11.620000 371.080000 54.820000 372.160000 ;
      RECT 4.860000 371.080000 9.655000 372.160000 ;
      RECT 0.000000 371.080000 3.060000 372.160000 ;
      RECT 0.000000 369.810000 550.160000 371.080000 ;
      RECT 0.000000 369.440000 548.960000 369.810000 ;
      RECT 544.900000 368.830000 548.960000 369.440000 ;
      RECT 544.900000 368.360000 550.160000 368.830000 ;
      RECT 508.620000 368.360000 543.100000 369.440000 ;
      RECT 463.620000 368.360000 506.820000 369.440000 ;
      RECT 418.620000 368.360000 461.820000 369.440000 ;
      RECT 373.620000 368.360000 416.820000 369.440000 ;
      RECT 328.620000 368.360000 371.820000 369.440000 ;
      RECT 283.620000 368.360000 326.820000 369.440000 ;
      RECT 238.620000 368.360000 281.820000 369.440000 ;
      RECT 193.620000 368.360000 236.820000 369.440000 ;
      RECT 148.620000 368.360000 191.820000 369.440000 ;
      RECT 103.620000 368.360000 146.820000 369.440000 ;
      RECT 58.620000 368.360000 101.820000 369.440000 ;
      RECT 13.620000 368.360000 56.820000 369.440000 ;
      RECT 7.060000 368.360000 11.820000 369.440000 ;
      RECT 0.000000 368.360000 5.260000 369.440000 ;
      RECT 0.000000 366.720000 550.160000 368.360000 ;
      RECT 547.100000 366.150000 550.160000 366.720000 ;
      RECT 547.100000 365.640000 548.960000 366.150000 ;
      RECT 506.620000 365.640000 545.300000 366.720000 ;
      RECT 461.620000 365.640000 504.820000 366.720000 ;
      RECT 416.620000 365.640000 459.820000 366.720000 ;
      RECT 371.620000 365.640000 414.820000 366.720000 ;
      RECT 326.620000 365.640000 369.820000 366.720000 ;
      RECT 281.620000 365.640000 324.820000 366.720000 ;
      RECT 236.620000 365.640000 279.820000 366.720000 ;
      RECT 191.620000 365.640000 234.820000 366.720000 ;
      RECT 146.620000 365.640000 189.820000 366.720000 ;
      RECT 101.620000 365.640000 144.820000 366.720000 ;
      RECT 56.620000 365.640000 99.820000 366.720000 ;
      RECT 11.620000 365.640000 54.820000 366.720000 ;
      RECT 4.860000 365.640000 9.655000 366.720000 ;
      RECT 0.000000 365.640000 3.060000 366.720000 ;
      RECT 0.000000 365.170000 548.960000 365.640000 ;
      RECT 0.000000 364.000000 550.160000 365.170000 ;
      RECT 544.900000 363.100000 550.160000 364.000000 ;
      RECT 544.900000 362.920000 548.960000 363.100000 ;
      RECT 508.620000 362.920000 543.100000 364.000000 ;
      RECT 463.620000 362.920000 506.820000 364.000000 ;
      RECT 418.620000 362.920000 461.820000 364.000000 ;
      RECT 373.620000 362.920000 416.820000 364.000000 ;
      RECT 328.620000 362.920000 371.820000 364.000000 ;
      RECT 283.620000 362.920000 326.820000 364.000000 ;
      RECT 238.620000 362.920000 281.820000 364.000000 ;
      RECT 193.620000 362.920000 236.820000 364.000000 ;
      RECT 148.620000 362.920000 191.820000 364.000000 ;
      RECT 103.620000 362.920000 146.820000 364.000000 ;
      RECT 58.620000 362.920000 101.820000 364.000000 ;
      RECT 13.620000 362.920000 56.820000 364.000000 ;
      RECT 7.060000 362.920000 11.820000 364.000000 ;
      RECT 0.000000 362.920000 5.260000 364.000000 ;
      RECT 0.000000 362.120000 548.960000 362.920000 ;
      RECT 0.000000 361.280000 550.160000 362.120000 ;
      RECT 547.100000 360.200000 550.160000 361.280000 ;
      RECT 506.620000 360.200000 545.300000 361.280000 ;
      RECT 461.620000 360.200000 504.820000 361.280000 ;
      RECT 416.620000 360.200000 459.820000 361.280000 ;
      RECT 371.620000 360.200000 414.820000 361.280000 ;
      RECT 326.620000 360.200000 369.820000 361.280000 ;
      RECT 281.620000 360.200000 324.820000 361.280000 ;
      RECT 236.620000 360.200000 279.820000 361.280000 ;
      RECT 191.620000 360.200000 234.820000 361.280000 ;
      RECT 146.620000 360.200000 189.820000 361.280000 ;
      RECT 101.620000 360.200000 144.820000 361.280000 ;
      RECT 56.620000 360.200000 99.820000 361.280000 ;
      RECT 11.620000 360.200000 54.820000 361.280000 ;
      RECT 4.860000 360.200000 9.655000 361.280000 ;
      RECT 0.000000 360.200000 3.060000 361.280000 ;
      RECT 0.000000 360.050000 550.160000 360.200000 ;
      RECT 0.000000 359.070000 548.960000 360.050000 ;
      RECT 0.000000 358.560000 550.160000 359.070000 ;
      RECT 544.900000 357.480000 550.160000 358.560000 ;
      RECT 508.620000 357.480000 543.100000 358.560000 ;
      RECT 463.620000 357.480000 506.820000 358.560000 ;
      RECT 418.620000 357.480000 461.820000 358.560000 ;
      RECT 373.620000 357.480000 416.820000 358.560000 ;
      RECT 328.620000 357.480000 371.820000 358.560000 ;
      RECT 283.620000 357.480000 326.820000 358.560000 ;
      RECT 238.620000 357.480000 281.820000 358.560000 ;
      RECT 193.620000 357.480000 236.820000 358.560000 ;
      RECT 148.620000 357.480000 191.820000 358.560000 ;
      RECT 103.620000 357.480000 146.820000 358.560000 ;
      RECT 58.620000 357.480000 101.820000 358.560000 ;
      RECT 13.620000 357.480000 56.820000 358.560000 ;
      RECT 7.060000 357.480000 11.820000 358.560000 ;
      RECT 0.000000 357.480000 5.260000 358.560000 ;
      RECT 0.000000 357.000000 550.160000 357.480000 ;
      RECT 0.000000 356.020000 548.960000 357.000000 ;
      RECT 0.000000 355.840000 550.160000 356.020000 ;
      RECT 547.100000 354.760000 550.160000 355.840000 ;
      RECT 506.620000 354.760000 545.300000 355.840000 ;
      RECT 461.620000 354.760000 504.820000 355.840000 ;
      RECT 416.620000 354.760000 459.820000 355.840000 ;
      RECT 371.620000 354.760000 414.820000 355.840000 ;
      RECT 326.620000 354.760000 369.820000 355.840000 ;
      RECT 281.620000 354.760000 324.820000 355.840000 ;
      RECT 236.620000 354.760000 279.820000 355.840000 ;
      RECT 191.620000 354.760000 234.820000 355.840000 ;
      RECT 146.620000 354.760000 189.820000 355.840000 ;
      RECT 101.620000 354.760000 144.820000 355.840000 ;
      RECT 56.620000 354.760000 99.820000 355.840000 ;
      RECT 11.620000 354.760000 54.820000 355.840000 ;
      RECT 4.860000 354.760000 9.655000 355.840000 ;
      RECT 0.000000 354.760000 3.060000 355.840000 ;
      RECT 0.000000 353.950000 550.160000 354.760000 ;
      RECT 0.000000 353.120000 548.960000 353.950000 ;
      RECT 544.900000 352.970000 548.960000 353.120000 ;
      RECT 544.900000 352.040000 550.160000 352.970000 ;
      RECT 508.620000 352.040000 543.100000 353.120000 ;
      RECT 463.620000 352.040000 506.820000 353.120000 ;
      RECT 418.620000 352.040000 461.820000 353.120000 ;
      RECT 373.620000 352.040000 416.820000 353.120000 ;
      RECT 328.620000 352.040000 371.820000 353.120000 ;
      RECT 283.620000 352.040000 326.820000 353.120000 ;
      RECT 238.620000 352.040000 281.820000 353.120000 ;
      RECT 193.620000 352.040000 236.820000 353.120000 ;
      RECT 148.620000 352.040000 191.820000 353.120000 ;
      RECT 103.620000 352.040000 146.820000 353.120000 ;
      RECT 58.620000 352.040000 101.820000 353.120000 ;
      RECT 13.620000 352.040000 56.820000 353.120000 ;
      RECT 7.060000 352.040000 11.820000 353.120000 ;
      RECT 0.000000 352.040000 5.260000 353.120000 ;
      RECT 0.000000 350.900000 550.160000 352.040000 ;
      RECT 0.000000 350.400000 548.960000 350.900000 ;
      RECT 547.100000 349.920000 548.960000 350.400000 ;
      RECT 547.100000 349.320000 550.160000 349.920000 ;
      RECT 506.620000 349.320000 545.300000 350.400000 ;
      RECT 461.620000 349.320000 504.820000 350.400000 ;
      RECT 416.620000 349.320000 459.820000 350.400000 ;
      RECT 371.620000 349.320000 414.820000 350.400000 ;
      RECT 326.620000 349.320000 369.820000 350.400000 ;
      RECT 281.620000 349.320000 324.820000 350.400000 ;
      RECT 236.620000 349.320000 279.820000 350.400000 ;
      RECT 191.620000 349.320000 234.820000 350.400000 ;
      RECT 146.620000 349.320000 189.820000 350.400000 ;
      RECT 101.620000 349.320000 144.820000 350.400000 ;
      RECT 56.620000 349.320000 99.820000 350.400000 ;
      RECT 11.620000 349.320000 54.820000 350.400000 ;
      RECT 4.860000 349.320000 9.655000 350.400000 ;
      RECT 0.000000 349.320000 3.060000 350.400000 ;
      RECT 0.000000 347.680000 550.160000 349.320000 ;
      RECT 544.900000 347.240000 550.160000 347.680000 ;
      RECT 544.900000 346.600000 548.960000 347.240000 ;
      RECT 508.620000 346.600000 543.100000 347.680000 ;
      RECT 463.620000 346.600000 506.820000 347.680000 ;
      RECT 418.620000 346.600000 461.820000 347.680000 ;
      RECT 373.620000 346.600000 416.820000 347.680000 ;
      RECT 328.620000 346.600000 371.820000 347.680000 ;
      RECT 283.620000 346.600000 326.820000 347.680000 ;
      RECT 238.620000 346.600000 281.820000 347.680000 ;
      RECT 193.620000 346.600000 236.820000 347.680000 ;
      RECT 148.620000 346.600000 191.820000 347.680000 ;
      RECT 103.620000 346.600000 146.820000 347.680000 ;
      RECT 58.620000 346.600000 101.820000 347.680000 ;
      RECT 13.620000 346.600000 56.820000 347.680000 ;
      RECT 7.060000 346.600000 11.820000 347.680000 ;
      RECT 0.000000 346.600000 5.260000 347.680000 ;
      RECT 0.000000 346.260000 548.960000 346.600000 ;
      RECT 0.000000 344.960000 550.160000 346.260000 ;
      RECT 547.100000 344.190000 550.160000 344.960000 ;
      RECT 547.100000 343.880000 548.960000 344.190000 ;
      RECT 506.620000 343.880000 545.300000 344.960000 ;
      RECT 461.620000 343.880000 504.820000 344.960000 ;
      RECT 416.620000 343.880000 459.820000 344.960000 ;
      RECT 371.620000 343.880000 414.820000 344.960000 ;
      RECT 326.620000 343.880000 369.820000 344.960000 ;
      RECT 281.620000 343.880000 324.820000 344.960000 ;
      RECT 236.620000 343.880000 279.820000 344.960000 ;
      RECT 191.620000 343.880000 234.820000 344.960000 ;
      RECT 146.620000 343.880000 189.820000 344.960000 ;
      RECT 101.620000 343.880000 144.820000 344.960000 ;
      RECT 56.620000 343.880000 99.820000 344.960000 ;
      RECT 11.620000 343.880000 54.820000 344.960000 ;
      RECT 4.860000 343.880000 9.655000 344.960000 ;
      RECT 0.000000 343.880000 3.060000 344.960000 ;
      RECT 0.000000 343.210000 548.960000 343.880000 ;
      RECT 0.000000 342.240000 550.160000 343.210000 ;
      RECT 544.900000 341.160000 550.160000 342.240000 ;
      RECT 508.620000 341.160000 543.100000 342.240000 ;
      RECT 463.620000 341.160000 506.820000 342.240000 ;
      RECT 418.620000 341.160000 461.820000 342.240000 ;
      RECT 373.620000 341.160000 416.820000 342.240000 ;
      RECT 328.620000 341.160000 371.820000 342.240000 ;
      RECT 283.620000 341.160000 326.820000 342.240000 ;
      RECT 238.620000 341.160000 281.820000 342.240000 ;
      RECT 193.620000 341.160000 236.820000 342.240000 ;
      RECT 148.620000 341.160000 191.820000 342.240000 ;
      RECT 103.620000 341.160000 146.820000 342.240000 ;
      RECT 58.620000 341.160000 101.820000 342.240000 ;
      RECT 13.620000 341.160000 56.820000 342.240000 ;
      RECT 7.060000 341.160000 11.820000 342.240000 ;
      RECT 0.000000 341.160000 5.260000 342.240000 ;
      RECT 0.000000 341.140000 550.160000 341.160000 ;
      RECT 0.000000 340.160000 548.960000 341.140000 ;
      RECT 0.000000 339.520000 550.160000 340.160000 ;
      RECT 547.100000 338.440000 550.160000 339.520000 ;
      RECT 506.620000 338.440000 545.300000 339.520000 ;
      RECT 461.620000 338.440000 504.820000 339.520000 ;
      RECT 416.620000 338.440000 459.820000 339.520000 ;
      RECT 371.620000 338.440000 414.820000 339.520000 ;
      RECT 326.620000 338.440000 369.820000 339.520000 ;
      RECT 281.620000 338.440000 324.820000 339.520000 ;
      RECT 236.620000 338.440000 279.820000 339.520000 ;
      RECT 191.620000 338.440000 234.820000 339.520000 ;
      RECT 146.620000 338.440000 189.820000 339.520000 ;
      RECT 101.620000 338.440000 144.820000 339.520000 ;
      RECT 56.620000 338.440000 99.820000 339.520000 ;
      RECT 11.620000 338.440000 54.820000 339.520000 ;
      RECT 4.860000 338.440000 9.655000 339.520000 ;
      RECT 0.000000 338.440000 3.060000 339.520000 ;
      RECT 0.000000 338.090000 550.160000 338.440000 ;
      RECT 0.000000 337.110000 548.960000 338.090000 ;
      RECT 0.000000 336.800000 550.160000 337.110000 ;
      RECT 544.900000 335.720000 550.160000 336.800000 ;
      RECT 508.620000 335.720000 543.100000 336.800000 ;
      RECT 463.620000 335.720000 506.820000 336.800000 ;
      RECT 418.620000 335.720000 461.820000 336.800000 ;
      RECT 373.620000 335.720000 416.820000 336.800000 ;
      RECT 328.620000 335.720000 371.820000 336.800000 ;
      RECT 283.620000 335.720000 326.820000 336.800000 ;
      RECT 238.620000 335.720000 281.820000 336.800000 ;
      RECT 193.620000 335.720000 236.820000 336.800000 ;
      RECT 148.620000 335.720000 191.820000 336.800000 ;
      RECT 103.620000 335.720000 146.820000 336.800000 ;
      RECT 58.620000 335.720000 101.820000 336.800000 ;
      RECT 13.620000 335.720000 56.820000 336.800000 ;
      RECT 7.060000 335.720000 11.820000 336.800000 ;
      RECT 0.000000 335.720000 5.260000 336.800000 ;
      RECT 0.000000 335.040000 550.160000 335.720000 ;
      RECT 0.000000 334.080000 548.960000 335.040000 ;
      RECT 547.100000 334.060000 548.960000 334.080000 ;
      RECT 547.100000 333.000000 550.160000 334.060000 ;
      RECT 506.620000 333.000000 545.300000 334.080000 ;
      RECT 461.620000 333.000000 504.820000 334.080000 ;
      RECT 416.620000 333.000000 459.820000 334.080000 ;
      RECT 371.620000 333.000000 414.820000 334.080000 ;
      RECT 326.620000 333.000000 369.820000 334.080000 ;
      RECT 281.620000 333.000000 324.820000 334.080000 ;
      RECT 236.620000 333.000000 279.820000 334.080000 ;
      RECT 191.620000 333.000000 234.820000 334.080000 ;
      RECT 146.620000 333.000000 189.820000 334.080000 ;
      RECT 101.620000 333.000000 144.820000 334.080000 ;
      RECT 56.620000 333.000000 99.820000 334.080000 ;
      RECT 11.620000 333.000000 54.820000 334.080000 ;
      RECT 4.860000 333.000000 9.655000 334.080000 ;
      RECT 0.000000 333.000000 3.060000 334.080000 ;
      RECT 0.000000 331.990000 550.160000 333.000000 ;
      RECT 0.000000 331.360000 548.960000 331.990000 ;
      RECT 544.900000 331.010000 548.960000 331.360000 ;
      RECT 544.900000 330.280000 550.160000 331.010000 ;
      RECT 508.620000 330.280000 543.100000 331.360000 ;
      RECT 463.620000 330.280000 506.820000 331.360000 ;
      RECT 418.620000 330.280000 461.820000 331.360000 ;
      RECT 373.620000 330.280000 416.820000 331.360000 ;
      RECT 328.620000 330.280000 371.820000 331.360000 ;
      RECT 283.620000 330.280000 326.820000 331.360000 ;
      RECT 238.620000 330.280000 281.820000 331.360000 ;
      RECT 193.620000 330.280000 236.820000 331.360000 ;
      RECT 148.620000 330.280000 191.820000 331.360000 ;
      RECT 103.620000 330.280000 146.820000 331.360000 ;
      RECT 58.620000 330.280000 101.820000 331.360000 ;
      RECT 13.620000 330.280000 56.820000 331.360000 ;
      RECT 7.060000 330.280000 11.820000 331.360000 ;
      RECT 0.000000 330.280000 5.260000 331.360000 ;
      RECT 0.000000 328.640000 550.160000 330.280000 ;
      RECT 547.100000 328.330000 550.160000 328.640000 ;
      RECT 547.100000 327.560000 548.960000 328.330000 ;
      RECT 506.620000 327.560000 545.300000 328.640000 ;
      RECT 461.620000 327.560000 504.820000 328.640000 ;
      RECT 416.620000 327.560000 459.820000 328.640000 ;
      RECT 371.620000 327.560000 414.820000 328.640000 ;
      RECT 326.620000 327.560000 369.820000 328.640000 ;
      RECT 281.620000 327.560000 324.820000 328.640000 ;
      RECT 236.620000 327.560000 279.820000 328.640000 ;
      RECT 191.620000 327.560000 234.820000 328.640000 ;
      RECT 146.620000 327.560000 189.820000 328.640000 ;
      RECT 101.620000 327.560000 144.820000 328.640000 ;
      RECT 56.620000 327.560000 99.820000 328.640000 ;
      RECT 11.620000 327.560000 54.820000 328.640000 ;
      RECT 4.860000 327.560000 9.655000 328.640000 ;
      RECT 0.000000 327.560000 3.060000 328.640000 ;
      RECT 0.000000 327.350000 548.960000 327.560000 ;
      RECT 0.000000 325.920000 550.160000 327.350000 ;
      RECT 544.900000 325.280000 550.160000 325.920000 ;
      RECT 544.900000 324.840000 548.960000 325.280000 ;
      RECT 508.620000 324.840000 543.100000 325.920000 ;
      RECT 463.620000 324.840000 506.820000 325.920000 ;
      RECT 418.620000 324.840000 461.820000 325.920000 ;
      RECT 373.620000 324.840000 416.820000 325.920000 ;
      RECT 328.620000 324.840000 371.820000 325.920000 ;
      RECT 283.620000 324.840000 326.820000 325.920000 ;
      RECT 238.620000 324.840000 281.820000 325.920000 ;
      RECT 193.620000 324.840000 236.820000 325.920000 ;
      RECT 148.620000 324.840000 191.820000 325.920000 ;
      RECT 103.620000 324.840000 146.820000 325.920000 ;
      RECT 58.620000 324.840000 101.820000 325.920000 ;
      RECT 13.620000 324.840000 56.820000 325.920000 ;
      RECT 7.060000 324.840000 11.820000 325.920000 ;
      RECT 0.000000 324.840000 5.260000 325.920000 ;
      RECT 0.000000 324.300000 548.960000 324.840000 ;
      RECT 0.000000 323.200000 550.160000 324.300000 ;
      RECT 547.100000 322.230000 550.160000 323.200000 ;
      RECT 547.100000 322.120000 548.960000 322.230000 ;
      RECT 506.620000 322.120000 545.300000 323.200000 ;
      RECT 461.620000 322.120000 504.820000 323.200000 ;
      RECT 416.620000 322.120000 459.820000 323.200000 ;
      RECT 371.620000 322.120000 414.820000 323.200000 ;
      RECT 326.620000 322.120000 369.820000 323.200000 ;
      RECT 281.620000 322.120000 324.820000 323.200000 ;
      RECT 236.620000 322.120000 279.820000 323.200000 ;
      RECT 191.620000 322.120000 234.820000 323.200000 ;
      RECT 146.620000 322.120000 189.820000 323.200000 ;
      RECT 101.620000 322.120000 144.820000 323.200000 ;
      RECT 56.620000 322.120000 99.820000 323.200000 ;
      RECT 11.620000 322.120000 54.820000 323.200000 ;
      RECT 4.860000 322.120000 9.655000 323.200000 ;
      RECT 0.000000 322.120000 3.060000 323.200000 ;
      RECT 0.000000 321.250000 548.960000 322.120000 ;
      RECT 0.000000 320.480000 550.160000 321.250000 ;
      RECT 544.900000 319.400000 550.160000 320.480000 ;
      RECT 508.620000 319.400000 543.100000 320.480000 ;
      RECT 463.620000 319.400000 506.820000 320.480000 ;
      RECT 418.620000 319.400000 461.820000 320.480000 ;
      RECT 373.620000 319.400000 416.820000 320.480000 ;
      RECT 328.620000 319.400000 371.820000 320.480000 ;
      RECT 283.620000 319.400000 326.820000 320.480000 ;
      RECT 238.620000 319.400000 281.820000 320.480000 ;
      RECT 193.620000 319.400000 236.820000 320.480000 ;
      RECT 148.620000 319.400000 191.820000 320.480000 ;
      RECT 103.620000 319.400000 146.820000 320.480000 ;
      RECT 58.620000 319.400000 101.820000 320.480000 ;
      RECT 13.620000 319.400000 56.820000 320.480000 ;
      RECT 7.060000 319.400000 11.820000 320.480000 ;
      RECT 0.000000 319.400000 5.260000 320.480000 ;
      RECT 0.000000 319.180000 550.160000 319.400000 ;
      RECT 0.000000 318.200000 548.960000 319.180000 ;
      RECT 0.000000 317.760000 550.160000 318.200000 ;
      RECT 547.100000 316.680000 550.160000 317.760000 ;
      RECT 506.620000 316.680000 545.300000 317.760000 ;
      RECT 461.620000 316.680000 504.820000 317.760000 ;
      RECT 416.620000 316.680000 459.820000 317.760000 ;
      RECT 371.620000 316.680000 414.820000 317.760000 ;
      RECT 326.620000 316.680000 369.820000 317.760000 ;
      RECT 281.620000 316.680000 324.820000 317.760000 ;
      RECT 236.620000 316.680000 279.820000 317.760000 ;
      RECT 191.620000 316.680000 234.820000 317.760000 ;
      RECT 146.620000 316.680000 189.820000 317.760000 ;
      RECT 101.620000 316.680000 144.820000 317.760000 ;
      RECT 56.620000 316.680000 99.820000 317.760000 ;
      RECT 11.620000 316.680000 54.820000 317.760000 ;
      RECT 4.860000 316.680000 9.655000 317.760000 ;
      RECT 0.000000 316.680000 3.060000 317.760000 ;
      RECT 0.000000 316.130000 550.160000 316.680000 ;
      RECT 0.000000 315.150000 548.960000 316.130000 ;
      RECT 0.000000 315.040000 550.160000 315.150000 ;
      RECT 544.900000 313.960000 550.160000 315.040000 ;
      RECT 508.620000 313.960000 543.100000 315.040000 ;
      RECT 463.620000 313.960000 506.820000 315.040000 ;
      RECT 418.620000 313.960000 461.820000 315.040000 ;
      RECT 373.620000 313.960000 416.820000 315.040000 ;
      RECT 328.620000 313.960000 371.820000 315.040000 ;
      RECT 283.620000 313.960000 326.820000 315.040000 ;
      RECT 238.620000 313.960000 281.820000 315.040000 ;
      RECT 193.620000 313.960000 236.820000 315.040000 ;
      RECT 148.620000 313.960000 191.820000 315.040000 ;
      RECT 103.620000 313.960000 146.820000 315.040000 ;
      RECT 58.620000 313.960000 101.820000 315.040000 ;
      RECT 13.620000 313.960000 56.820000 315.040000 ;
      RECT 7.060000 313.960000 11.820000 315.040000 ;
      RECT 0.000000 313.960000 5.260000 315.040000 ;
      RECT 0.000000 313.080000 550.160000 313.960000 ;
      RECT 0.000000 312.320000 548.960000 313.080000 ;
      RECT 547.100000 312.100000 548.960000 312.320000 ;
      RECT 547.100000 311.240000 550.160000 312.100000 ;
      RECT 506.620000 311.240000 545.300000 312.320000 ;
      RECT 461.620000 311.240000 504.820000 312.320000 ;
      RECT 416.620000 311.240000 459.820000 312.320000 ;
      RECT 371.620000 311.240000 414.820000 312.320000 ;
      RECT 326.620000 311.240000 369.820000 312.320000 ;
      RECT 281.620000 311.240000 324.820000 312.320000 ;
      RECT 236.620000 311.240000 279.820000 312.320000 ;
      RECT 191.620000 311.240000 234.820000 312.320000 ;
      RECT 146.620000 311.240000 189.820000 312.320000 ;
      RECT 101.620000 311.240000 144.820000 312.320000 ;
      RECT 56.620000 311.240000 99.820000 312.320000 ;
      RECT 11.620000 311.240000 54.820000 312.320000 ;
      RECT 4.860000 311.240000 9.655000 312.320000 ;
      RECT 0.000000 311.240000 3.060000 312.320000 ;
      RECT 0.000000 309.600000 550.160000 311.240000 ;
      RECT 544.900000 309.420000 550.160000 309.600000 ;
      RECT 544.900000 308.520000 548.960000 309.420000 ;
      RECT 508.620000 308.520000 543.100000 309.600000 ;
      RECT 463.620000 308.520000 506.820000 309.600000 ;
      RECT 418.620000 308.520000 461.820000 309.600000 ;
      RECT 373.620000 308.520000 416.820000 309.600000 ;
      RECT 328.620000 308.520000 371.820000 309.600000 ;
      RECT 283.620000 308.520000 326.820000 309.600000 ;
      RECT 238.620000 308.520000 281.820000 309.600000 ;
      RECT 193.620000 308.520000 236.820000 309.600000 ;
      RECT 148.620000 308.520000 191.820000 309.600000 ;
      RECT 103.620000 308.520000 146.820000 309.600000 ;
      RECT 58.620000 308.520000 101.820000 309.600000 ;
      RECT 13.620000 308.520000 56.820000 309.600000 ;
      RECT 7.060000 308.520000 11.820000 309.600000 ;
      RECT 0.000000 308.520000 5.260000 309.600000 ;
      RECT 0.000000 308.440000 548.960000 308.520000 ;
      RECT 0.000000 306.880000 550.160000 308.440000 ;
      RECT 547.100000 306.370000 550.160000 306.880000 ;
      RECT 547.100000 305.800000 548.960000 306.370000 ;
      RECT 506.620000 305.800000 545.300000 306.880000 ;
      RECT 461.620000 305.800000 504.820000 306.880000 ;
      RECT 416.620000 305.800000 459.820000 306.880000 ;
      RECT 371.620000 305.800000 414.820000 306.880000 ;
      RECT 326.620000 305.800000 369.820000 306.880000 ;
      RECT 281.620000 305.800000 324.820000 306.880000 ;
      RECT 236.620000 305.800000 279.820000 306.880000 ;
      RECT 191.620000 305.800000 234.820000 306.880000 ;
      RECT 146.620000 305.800000 189.820000 306.880000 ;
      RECT 101.620000 305.800000 144.820000 306.880000 ;
      RECT 56.620000 305.800000 99.820000 306.880000 ;
      RECT 11.620000 305.800000 54.820000 306.880000 ;
      RECT 4.860000 305.800000 9.655000 306.880000 ;
      RECT 0.000000 305.800000 3.060000 306.880000 ;
      RECT 0.000000 305.390000 548.960000 305.800000 ;
      RECT 0.000000 304.160000 550.160000 305.390000 ;
      RECT 544.900000 303.320000 550.160000 304.160000 ;
      RECT 544.900000 303.080000 548.960000 303.320000 ;
      RECT 508.620000 303.080000 543.100000 304.160000 ;
      RECT 463.620000 303.080000 506.820000 304.160000 ;
      RECT 418.620000 303.080000 461.820000 304.160000 ;
      RECT 373.620000 303.080000 416.820000 304.160000 ;
      RECT 328.620000 303.080000 371.820000 304.160000 ;
      RECT 283.620000 303.080000 326.820000 304.160000 ;
      RECT 238.620000 303.080000 281.820000 304.160000 ;
      RECT 193.620000 303.080000 236.820000 304.160000 ;
      RECT 148.620000 303.080000 191.820000 304.160000 ;
      RECT 103.620000 303.080000 146.820000 304.160000 ;
      RECT 58.620000 303.080000 101.820000 304.160000 ;
      RECT 13.620000 303.080000 56.820000 304.160000 ;
      RECT 7.060000 303.080000 11.820000 304.160000 ;
      RECT 0.000000 303.080000 5.260000 304.160000 ;
      RECT 0.000000 302.340000 548.960000 303.080000 ;
      RECT 0.000000 301.440000 550.160000 302.340000 ;
      RECT 547.100000 300.360000 550.160000 301.440000 ;
      RECT 506.620000 300.360000 545.300000 301.440000 ;
      RECT 461.620000 300.360000 504.820000 301.440000 ;
      RECT 416.620000 300.360000 459.820000 301.440000 ;
      RECT 371.620000 300.360000 414.820000 301.440000 ;
      RECT 326.620000 300.360000 369.820000 301.440000 ;
      RECT 281.620000 300.360000 324.820000 301.440000 ;
      RECT 236.620000 300.360000 279.820000 301.440000 ;
      RECT 191.620000 300.360000 234.820000 301.440000 ;
      RECT 146.620000 300.360000 189.820000 301.440000 ;
      RECT 101.620000 300.360000 144.820000 301.440000 ;
      RECT 56.620000 300.360000 99.820000 301.440000 ;
      RECT 11.620000 300.360000 54.820000 301.440000 ;
      RECT 4.860000 300.360000 9.655000 301.440000 ;
      RECT 0.000000 300.360000 3.060000 301.440000 ;
      RECT 0.000000 300.270000 550.160000 300.360000 ;
      RECT 0.000000 299.290000 548.960000 300.270000 ;
      RECT 0.000000 298.720000 550.160000 299.290000 ;
      RECT 544.900000 297.640000 550.160000 298.720000 ;
      RECT 508.620000 297.640000 543.100000 298.720000 ;
      RECT 463.620000 297.640000 506.820000 298.720000 ;
      RECT 418.620000 297.640000 461.820000 298.720000 ;
      RECT 373.620000 297.640000 416.820000 298.720000 ;
      RECT 328.620000 297.640000 371.820000 298.720000 ;
      RECT 283.620000 297.640000 326.820000 298.720000 ;
      RECT 238.620000 297.640000 281.820000 298.720000 ;
      RECT 193.620000 297.640000 236.820000 298.720000 ;
      RECT 148.620000 297.640000 191.820000 298.720000 ;
      RECT 103.620000 297.640000 146.820000 298.720000 ;
      RECT 58.620000 297.640000 101.820000 298.720000 ;
      RECT 13.620000 297.640000 56.820000 298.720000 ;
      RECT 7.060000 297.640000 11.820000 298.720000 ;
      RECT 0.000000 297.640000 5.260000 298.720000 ;
      RECT 0.000000 297.220000 550.160000 297.640000 ;
      RECT 0.000000 296.240000 548.960000 297.220000 ;
      RECT 0.000000 296.000000 550.160000 296.240000 ;
      RECT 547.100000 294.920000 550.160000 296.000000 ;
      RECT 506.620000 294.920000 545.300000 296.000000 ;
      RECT 461.620000 294.920000 504.820000 296.000000 ;
      RECT 416.620000 294.920000 459.820000 296.000000 ;
      RECT 371.620000 294.920000 414.820000 296.000000 ;
      RECT 326.620000 294.920000 369.820000 296.000000 ;
      RECT 281.620000 294.920000 324.820000 296.000000 ;
      RECT 236.620000 294.920000 279.820000 296.000000 ;
      RECT 191.620000 294.920000 234.820000 296.000000 ;
      RECT 146.620000 294.920000 189.820000 296.000000 ;
      RECT 101.620000 294.920000 144.820000 296.000000 ;
      RECT 56.620000 294.920000 99.820000 296.000000 ;
      RECT 11.620000 294.920000 54.820000 296.000000 ;
      RECT 4.860000 294.920000 9.655000 296.000000 ;
      RECT 0.000000 294.920000 3.060000 296.000000 ;
      RECT 0.000000 294.170000 550.160000 294.920000 ;
      RECT 0.000000 293.280000 548.960000 294.170000 ;
      RECT 544.900000 293.190000 548.960000 293.280000 ;
      RECT 544.900000 292.200000 550.160000 293.190000 ;
      RECT 508.620000 292.200000 543.100000 293.280000 ;
      RECT 463.620000 292.200000 506.820000 293.280000 ;
      RECT 418.620000 292.200000 461.820000 293.280000 ;
      RECT 373.620000 292.200000 416.820000 293.280000 ;
      RECT 328.620000 292.200000 371.820000 293.280000 ;
      RECT 283.620000 292.200000 326.820000 293.280000 ;
      RECT 238.620000 292.200000 281.820000 293.280000 ;
      RECT 193.620000 292.200000 236.820000 293.280000 ;
      RECT 148.620000 292.200000 191.820000 293.280000 ;
      RECT 103.620000 292.200000 146.820000 293.280000 ;
      RECT 58.620000 292.200000 101.820000 293.280000 ;
      RECT 13.620000 292.200000 56.820000 293.280000 ;
      RECT 7.060000 292.200000 11.820000 293.280000 ;
      RECT 0.000000 292.200000 5.260000 293.280000 ;
      RECT 0.000000 290.560000 550.160000 292.200000 ;
      RECT 547.100000 290.510000 550.160000 290.560000 ;
      RECT 547.100000 289.530000 548.960000 290.510000 ;
      RECT 547.100000 289.480000 550.160000 289.530000 ;
      RECT 506.620000 289.480000 545.300000 290.560000 ;
      RECT 461.620000 289.480000 504.820000 290.560000 ;
      RECT 416.620000 289.480000 459.820000 290.560000 ;
      RECT 371.620000 289.480000 414.820000 290.560000 ;
      RECT 326.620000 289.480000 369.820000 290.560000 ;
      RECT 281.620000 289.480000 324.820000 290.560000 ;
      RECT 236.620000 289.480000 279.820000 290.560000 ;
      RECT 191.620000 289.480000 234.820000 290.560000 ;
      RECT 146.620000 289.480000 189.820000 290.560000 ;
      RECT 101.620000 289.480000 144.820000 290.560000 ;
      RECT 56.620000 289.480000 99.820000 290.560000 ;
      RECT 11.620000 289.480000 54.820000 290.560000 ;
      RECT 4.860000 289.480000 9.655000 290.560000 ;
      RECT 0.000000 289.480000 3.060000 290.560000 ;
      RECT 0.000000 287.840000 550.160000 289.480000 ;
      RECT 544.900000 287.460000 550.160000 287.840000 ;
      RECT 544.900000 286.760000 548.960000 287.460000 ;
      RECT 508.620000 286.760000 543.100000 287.840000 ;
      RECT 463.620000 286.760000 506.820000 287.840000 ;
      RECT 418.620000 286.760000 461.820000 287.840000 ;
      RECT 373.620000 286.760000 416.820000 287.840000 ;
      RECT 328.620000 286.760000 371.820000 287.840000 ;
      RECT 283.620000 286.760000 326.820000 287.840000 ;
      RECT 238.620000 286.760000 281.820000 287.840000 ;
      RECT 193.620000 286.760000 236.820000 287.840000 ;
      RECT 148.620000 286.760000 191.820000 287.840000 ;
      RECT 103.620000 286.760000 146.820000 287.840000 ;
      RECT 58.620000 286.760000 101.820000 287.840000 ;
      RECT 13.620000 286.760000 56.820000 287.840000 ;
      RECT 7.060000 286.760000 11.820000 287.840000 ;
      RECT 0.000000 286.760000 5.260000 287.840000 ;
      RECT 0.000000 286.480000 548.960000 286.760000 ;
      RECT 0.000000 285.120000 550.160000 286.480000 ;
      RECT 547.100000 284.410000 550.160000 285.120000 ;
      RECT 547.100000 284.040000 548.960000 284.410000 ;
      RECT 506.620000 284.040000 545.300000 285.120000 ;
      RECT 461.620000 284.040000 504.820000 285.120000 ;
      RECT 416.620000 284.040000 459.820000 285.120000 ;
      RECT 371.620000 284.040000 414.820000 285.120000 ;
      RECT 326.620000 284.040000 369.820000 285.120000 ;
      RECT 281.620000 284.040000 324.820000 285.120000 ;
      RECT 236.620000 284.040000 279.820000 285.120000 ;
      RECT 191.620000 284.040000 234.820000 285.120000 ;
      RECT 146.620000 284.040000 189.820000 285.120000 ;
      RECT 101.620000 284.040000 144.820000 285.120000 ;
      RECT 56.620000 284.040000 99.820000 285.120000 ;
      RECT 11.620000 284.040000 54.820000 285.120000 ;
      RECT 4.860000 284.040000 9.655000 285.120000 ;
      RECT 0.000000 284.040000 3.060000 285.120000 ;
      RECT 0.000000 283.430000 548.960000 284.040000 ;
      RECT 0.000000 282.400000 550.160000 283.430000 ;
      RECT 544.900000 281.360000 550.160000 282.400000 ;
      RECT 544.900000 281.320000 548.960000 281.360000 ;
      RECT 508.620000 281.320000 543.100000 282.400000 ;
      RECT 463.620000 281.320000 506.820000 282.400000 ;
      RECT 418.620000 281.320000 461.820000 282.400000 ;
      RECT 373.620000 281.320000 416.820000 282.400000 ;
      RECT 328.620000 281.320000 371.820000 282.400000 ;
      RECT 283.620000 281.320000 326.820000 282.400000 ;
      RECT 238.620000 281.320000 281.820000 282.400000 ;
      RECT 193.620000 281.320000 236.820000 282.400000 ;
      RECT 148.620000 281.320000 191.820000 282.400000 ;
      RECT 103.620000 281.320000 146.820000 282.400000 ;
      RECT 58.620000 281.320000 101.820000 282.400000 ;
      RECT 13.620000 281.320000 56.820000 282.400000 ;
      RECT 7.060000 281.320000 11.820000 282.400000 ;
      RECT 0.000000 281.320000 5.260000 282.400000 ;
      RECT 0.000000 280.380000 548.960000 281.320000 ;
      RECT 0.000000 279.680000 550.160000 280.380000 ;
      RECT 547.100000 278.600000 550.160000 279.680000 ;
      RECT 506.620000 278.600000 545.300000 279.680000 ;
      RECT 461.620000 278.600000 504.820000 279.680000 ;
      RECT 416.620000 278.600000 459.820000 279.680000 ;
      RECT 371.620000 278.600000 414.820000 279.680000 ;
      RECT 326.620000 278.600000 369.820000 279.680000 ;
      RECT 281.620000 278.600000 324.820000 279.680000 ;
      RECT 236.620000 278.600000 279.820000 279.680000 ;
      RECT 191.620000 278.600000 234.820000 279.680000 ;
      RECT 146.620000 278.600000 189.820000 279.680000 ;
      RECT 101.620000 278.600000 144.820000 279.680000 ;
      RECT 56.620000 278.600000 99.820000 279.680000 ;
      RECT 11.620000 278.600000 54.820000 279.680000 ;
      RECT 4.860000 278.600000 9.655000 279.680000 ;
      RECT 0.000000 278.600000 3.060000 279.680000 ;
      RECT 0.000000 278.310000 550.160000 278.600000 ;
      RECT 0.000000 277.330000 548.960000 278.310000 ;
      RECT 0.000000 276.960000 550.160000 277.330000 ;
      RECT 544.900000 275.880000 550.160000 276.960000 ;
      RECT 508.620000 275.880000 543.100000 276.960000 ;
      RECT 463.620000 275.880000 506.820000 276.960000 ;
      RECT 418.620000 275.880000 461.820000 276.960000 ;
      RECT 373.620000 275.880000 416.820000 276.960000 ;
      RECT 328.620000 275.880000 371.820000 276.960000 ;
      RECT 283.620000 275.880000 326.820000 276.960000 ;
      RECT 238.620000 275.880000 281.820000 276.960000 ;
      RECT 193.620000 275.880000 236.820000 276.960000 ;
      RECT 148.620000 275.880000 191.820000 276.960000 ;
      RECT 103.620000 275.880000 146.820000 276.960000 ;
      RECT 58.620000 275.880000 101.820000 276.960000 ;
      RECT 13.620000 275.880000 56.820000 276.960000 ;
      RECT 7.060000 275.880000 11.820000 276.960000 ;
      RECT 0.000000 275.880000 5.260000 276.960000 ;
      RECT 0.000000 275.260000 550.160000 275.880000 ;
      RECT 0.000000 274.280000 548.960000 275.260000 ;
      RECT 0.000000 274.240000 550.160000 274.280000 ;
      RECT 547.100000 273.160000 550.160000 274.240000 ;
      RECT 506.620000 273.160000 545.300000 274.240000 ;
      RECT 461.620000 273.160000 504.820000 274.240000 ;
      RECT 416.620000 273.160000 459.820000 274.240000 ;
      RECT 371.620000 273.160000 414.820000 274.240000 ;
      RECT 326.620000 273.160000 369.820000 274.240000 ;
      RECT 281.620000 273.160000 324.820000 274.240000 ;
      RECT 236.620000 273.160000 279.820000 274.240000 ;
      RECT 191.620000 273.160000 234.820000 274.240000 ;
      RECT 146.620000 273.160000 189.820000 274.240000 ;
      RECT 101.620000 273.160000 144.820000 274.240000 ;
      RECT 56.620000 273.160000 99.820000 274.240000 ;
      RECT 11.620000 273.160000 54.820000 274.240000 ;
      RECT 4.860000 273.160000 9.655000 274.240000 ;
      RECT 0.000000 273.160000 3.060000 274.240000 ;
      RECT 0.000000 271.600000 550.160000 273.160000 ;
      RECT 0.000000 271.520000 548.960000 271.600000 ;
      RECT 544.900000 270.620000 548.960000 271.520000 ;
      RECT 544.900000 270.440000 550.160000 270.620000 ;
      RECT 508.620000 270.440000 543.100000 271.520000 ;
      RECT 463.620000 270.440000 506.820000 271.520000 ;
      RECT 418.620000 270.440000 461.820000 271.520000 ;
      RECT 373.620000 270.440000 416.820000 271.520000 ;
      RECT 328.620000 270.440000 371.820000 271.520000 ;
      RECT 283.620000 270.440000 326.820000 271.520000 ;
      RECT 238.620000 270.440000 281.820000 271.520000 ;
      RECT 193.620000 270.440000 236.820000 271.520000 ;
      RECT 148.620000 270.440000 191.820000 271.520000 ;
      RECT 103.620000 270.440000 146.820000 271.520000 ;
      RECT 58.620000 270.440000 101.820000 271.520000 ;
      RECT 13.620000 270.440000 56.820000 271.520000 ;
      RECT 7.060000 270.440000 11.820000 271.520000 ;
      RECT 0.000000 270.440000 5.260000 271.520000 ;
      RECT 0.000000 268.800000 550.160000 270.440000 ;
      RECT 547.100000 268.550000 550.160000 268.800000 ;
      RECT 547.100000 267.720000 548.960000 268.550000 ;
      RECT 506.620000 267.720000 545.300000 268.800000 ;
      RECT 461.620000 267.720000 504.820000 268.800000 ;
      RECT 416.620000 267.720000 459.820000 268.800000 ;
      RECT 371.620000 267.720000 414.820000 268.800000 ;
      RECT 326.620000 267.720000 369.820000 268.800000 ;
      RECT 281.620000 267.720000 324.820000 268.800000 ;
      RECT 236.620000 267.720000 279.820000 268.800000 ;
      RECT 191.620000 267.720000 234.820000 268.800000 ;
      RECT 146.620000 267.720000 189.820000 268.800000 ;
      RECT 101.620000 267.720000 144.820000 268.800000 ;
      RECT 56.620000 267.720000 99.820000 268.800000 ;
      RECT 11.620000 267.720000 54.820000 268.800000 ;
      RECT 4.860000 267.720000 9.655000 268.800000 ;
      RECT 0.000000 267.720000 3.060000 268.800000 ;
      RECT 0.000000 267.570000 548.960000 267.720000 ;
      RECT 0.000000 266.080000 550.160000 267.570000 ;
      RECT 544.900000 265.500000 550.160000 266.080000 ;
      RECT 544.900000 265.000000 548.960000 265.500000 ;
      RECT 508.620000 265.000000 543.100000 266.080000 ;
      RECT 463.620000 265.000000 506.820000 266.080000 ;
      RECT 418.620000 265.000000 461.820000 266.080000 ;
      RECT 373.620000 265.000000 416.820000 266.080000 ;
      RECT 328.620000 265.000000 371.820000 266.080000 ;
      RECT 283.620000 265.000000 326.820000 266.080000 ;
      RECT 238.620000 265.000000 281.820000 266.080000 ;
      RECT 193.620000 265.000000 236.820000 266.080000 ;
      RECT 148.620000 265.000000 191.820000 266.080000 ;
      RECT 103.620000 265.000000 146.820000 266.080000 ;
      RECT 58.620000 265.000000 101.820000 266.080000 ;
      RECT 13.620000 265.000000 56.820000 266.080000 ;
      RECT 7.060000 265.000000 11.820000 266.080000 ;
      RECT 0.000000 265.000000 5.260000 266.080000 ;
      RECT 0.000000 264.520000 548.960000 265.000000 ;
      RECT 0.000000 263.360000 550.160000 264.520000 ;
      RECT 547.100000 262.450000 550.160000 263.360000 ;
      RECT 547.100000 262.280000 548.960000 262.450000 ;
      RECT 506.620000 262.280000 545.300000 263.360000 ;
      RECT 461.620000 262.280000 504.820000 263.360000 ;
      RECT 416.620000 262.280000 459.820000 263.360000 ;
      RECT 371.620000 262.280000 414.820000 263.360000 ;
      RECT 326.620000 262.280000 369.820000 263.360000 ;
      RECT 281.620000 262.280000 324.820000 263.360000 ;
      RECT 236.620000 262.280000 279.820000 263.360000 ;
      RECT 191.620000 262.280000 234.820000 263.360000 ;
      RECT 146.620000 262.280000 189.820000 263.360000 ;
      RECT 101.620000 262.280000 144.820000 263.360000 ;
      RECT 56.620000 262.280000 99.820000 263.360000 ;
      RECT 11.620000 262.280000 54.820000 263.360000 ;
      RECT 4.860000 262.280000 9.655000 263.360000 ;
      RECT 0.000000 262.280000 3.060000 263.360000 ;
      RECT 0.000000 261.470000 548.960000 262.280000 ;
      RECT 0.000000 260.640000 550.160000 261.470000 ;
      RECT 544.900000 259.560000 550.160000 260.640000 ;
      RECT 508.620000 259.560000 543.100000 260.640000 ;
      RECT 463.620000 259.560000 506.820000 260.640000 ;
      RECT 418.620000 259.560000 461.820000 260.640000 ;
      RECT 373.620000 259.560000 416.820000 260.640000 ;
      RECT 328.620000 259.560000 371.820000 260.640000 ;
      RECT 283.620000 259.560000 326.820000 260.640000 ;
      RECT 238.620000 259.560000 281.820000 260.640000 ;
      RECT 193.620000 259.560000 236.820000 260.640000 ;
      RECT 148.620000 259.560000 191.820000 260.640000 ;
      RECT 103.620000 259.560000 146.820000 260.640000 ;
      RECT 58.620000 259.560000 101.820000 260.640000 ;
      RECT 13.620000 259.560000 56.820000 260.640000 ;
      RECT 7.060000 259.560000 11.820000 260.640000 ;
      RECT 0.000000 259.560000 5.260000 260.640000 ;
      RECT 0.000000 259.400000 550.160000 259.560000 ;
      RECT 0.000000 258.420000 548.960000 259.400000 ;
      RECT 0.000000 257.920000 550.160000 258.420000 ;
      RECT 547.100000 256.840000 550.160000 257.920000 ;
      RECT 506.620000 256.840000 545.300000 257.920000 ;
      RECT 461.620000 256.840000 504.820000 257.920000 ;
      RECT 416.620000 256.840000 459.820000 257.920000 ;
      RECT 371.620000 256.840000 414.820000 257.920000 ;
      RECT 326.620000 256.840000 369.820000 257.920000 ;
      RECT 281.620000 256.840000 324.820000 257.920000 ;
      RECT 236.620000 256.840000 279.820000 257.920000 ;
      RECT 191.620000 256.840000 234.820000 257.920000 ;
      RECT 146.620000 256.840000 189.820000 257.920000 ;
      RECT 101.620000 256.840000 144.820000 257.920000 ;
      RECT 56.620000 256.840000 99.820000 257.920000 ;
      RECT 11.620000 256.840000 54.820000 257.920000 ;
      RECT 4.860000 256.840000 9.655000 257.920000 ;
      RECT 0.000000 256.840000 3.060000 257.920000 ;
      RECT 0.000000 256.350000 550.160000 256.840000 ;
      RECT 0.000000 255.370000 548.960000 256.350000 ;
      RECT 0.000000 255.200000 550.160000 255.370000 ;
      RECT 544.900000 254.120000 550.160000 255.200000 ;
      RECT 508.620000 254.120000 543.100000 255.200000 ;
      RECT 463.620000 254.120000 506.820000 255.200000 ;
      RECT 418.620000 254.120000 461.820000 255.200000 ;
      RECT 373.620000 254.120000 416.820000 255.200000 ;
      RECT 328.620000 254.120000 371.820000 255.200000 ;
      RECT 283.620000 254.120000 326.820000 255.200000 ;
      RECT 238.620000 254.120000 281.820000 255.200000 ;
      RECT 193.620000 254.120000 236.820000 255.200000 ;
      RECT 148.620000 254.120000 191.820000 255.200000 ;
      RECT 103.620000 254.120000 146.820000 255.200000 ;
      RECT 58.620000 254.120000 101.820000 255.200000 ;
      RECT 13.620000 254.120000 56.820000 255.200000 ;
      RECT 7.060000 254.120000 11.820000 255.200000 ;
      RECT 0.000000 254.120000 5.260000 255.200000 ;
      RECT 0.000000 252.690000 550.160000 254.120000 ;
      RECT 0.000000 252.480000 548.960000 252.690000 ;
      RECT 547.100000 251.710000 548.960000 252.480000 ;
      RECT 547.100000 251.400000 550.160000 251.710000 ;
      RECT 506.620000 251.400000 545.300000 252.480000 ;
      RECT 461.620000 251.400000 504.820000 252.480000 ;
      RECT 416.620000 251.400000 459.820000 252.480000 ;
      RECT 371.620000 251.400000 414.820000 252.480000 ;
      RECT 326.620000 251.400000 369.820000 252.480000 ;
      RECT 281.620000 251.400000 324.820000 252.480000 ;
      RECT 236.620000 251.400000 279.820000 252.480000 ;
      RECT 191.620000 251.400000 234.820000 252.480000 ;
      RECT 146.620000 251.400000 189.820000 252.480000 ;
      RECT 101.620000 251.400000 144.820000 252.480000 ;
      RECT 56.620000 251.400000 99.820000 252.480000 ;
      RECT 11.620000 251.400000 54.820000 252.480000 ;
      RECT 4.860000 251.400000 9.655000 252.480000 ;
      RECT 0.000000 251.400000 3.060000 252.480000 ;
      RECT 0.000000 249.760000 550.160000 251.400000 ;
      RECT 544.900000 249.640000 550.160000 249.760000 ;
      RECT 544.900000 248.680000 548.960000 249.640000 ;
      RECT 508.620000 248.680000 543.100000 249.760000 ;
      RECT 463.620000 248.680000 506.820000 249.760000 ;
      RECT 418.620000 248.680000 461.820000 249.760000 ;
      RECT 373.620000 248.680000 416.820000 249.760000 ;
      RECT 328.620000 248.680000 371.820000 249.760000 ;
      RECT 283.620000 248.680000 326.820000 249.760000 ;
      RECT 238.620000 248.680000 281.820000 249.760000 ;
      RECT 193.620000 248.680000 236.820000 249.760000 ;
      RECT 148.620000 248.680000 191.820000 249.760000 ;
      RECT 103.620000 248.680000 146.820000 249.760000 ;
      RECT 58.620000 248.680000 101.820000 249.760000 ;
      RECT 13.620000 248.680000 56.820000 249.760000 ;
      RECT 7.060000 248.680000 11.820000 249.760000 ;
      RECT 0.000000 248.680000 5.260000 249.760000 ;
      RECT 0.000000 248.660000 548.960000 248.680000 ;
      RECT 0.000000 247.040000 550.160000 248.660000 ;
      RECT 547.100000 246.590000 550.160000 247.040000 ;
      RECT 547.100000 245.960000 548.960000 246.590000 ;
      RECT 506.620000 245.960000 545.300000 247.040000 ;
      RECT 461.620000 245.960000 504.820000 247.040000 ;
      RECT 416.620000 245.960000 459.820000 247.040000 ;
      RECT 371.620000 245.960000 414.820000 247.040000 ;
      RECT 326.620000 245.960000 369.820000 247.040000 ;
      RECT 281.620000 245.960000 324.820000 247.040000 ;
      RECT 236.620000 245.960000 279.820000 247.040000 ;
      RECT 191.620000 245.960000 234.820000 247.040000 ;
      RECT 146.620000 245.960000 189.820000 247.040000 ;
      RECT 101.620000 245.960000 144.820000 247.040000 ;
      RECT 56.620000 245.960000 99.820000 247.040000 ;
      RECT 11.620000 245.960000 54.820000 247.040000 ;
      RECT 4.860000 245.960000 9.655000 247.040000 ;
      RECT 0.000000 245.960000 3.060000 247.040000 ;
      RECT 0.000000 245.610000 548.960000 245.960000 ;
      RECT 0.000000 244.320000 550.160000 245.610000 ;
      RECT 544.900000 243.540000 550.160000 244.320000 ;
      RECT 544.900000 243.240000 548.960000 243.540000 ;
      RECT 508.620000 243.240000 543.100000 244.320000 ;
      RECT 463.620000 243.240000 506.820000 244.320000 ;
      RECT 418.620000 243.240000 461.820000 244.320000 ;
      RECT 373.620000 243.240000 416.820000 244.320000 ;
      RECT 328.620000 243.240000 371.820000 244.320000 ;
      RECT 283.620000 243.240000 326.820000 244.320000 ;
      RECT 238.620000 243.240000 281.820000 244.320000 ;
      RECT 193.620000 243.240000 236.820000 244.320000 ;
      RECT 148.620000 243.240000 191.820000 244.320000 ;
      RECT 103.620000 243.240000 146.820000 244.320000 ;
      RECT 58.620000 243.240000 101.820000 244.320000 ;
      RECT 13.620000 243.240000 56.820000 244.320000 ;
      RECT 7.060000 243.240000 11.820000 244.320000 ;
      RECT 0.000000 243.240000 5.260000 244.320000 ;
      RECT 0.000000 242.560000 548.960000 243.240000 ;
      RECT 0.000000 241.600000 550.160000 242.560000 ;
      RECT 547.100000 240.520000 550.160000 241.600000 ;
      RECT 506.620000 240.520000 545.300000 241.600000 ;
      RECT 461.620000 240.520000 504.820000 241.600000 ;
      RECT 416.620000 240.520000 459.820000 241.600000 ;
      RECT 371.620000 240.520000 414.820000 241.600000 ;
      RECT 326.620000 240.520000 369.820000 241.600000 ;
      RECT 281.620000 240.520000 324.820000 241.600000 ;
      RECT 236.620000 240.520000 279.820000 241.600000 ;
      RECT 191.620000 240.520000 234.820000 241.600000 ;
      RECT 146.620000 240.520000 189.820000 241.600000 ;
      RECT 101.620000 240.520000 144.820000 241.600000 ;
      RECT 56.620000 240.520000 99.820000 241.600000 ;
      RECT 11.620000 240.520000 54.820000 241.600000 ;
      RECT 4.860000 240.520000 9.655000 241.600000 ;
      RECT 0.000000 240.520000 3.060000 241.600000 ;
      RECT 0.000000 240.490000 550.160000 240.520000 ;
      RECT 0.000000 239.510000 548.960000 240.490000 ;
      RECT 0.000000 238.880000 550.160000 239.510000 ;
      RECT 544.900000 237.800000 550.160000 238.880000 ;
      RECT 508.620000 237.800000 543.100000 238.880000 ;
      RECT 463.620000 237.800000 506.820000 238.880000 ;
      RECT 418.620000 237.800000 461.820000 238.880000 ;
      RECT 373.620000 237.800000 416.820000 238.880000 ;
      RECT 328.620000 237.800000 371.820000 238.880000 ;
      RECT 283.620000 237.800000 326.820000 238.880000 ;
      RECT 238.620000 237.800000 281.820000 238.880000 ;
      RECT 193.620000 237.800000 236.820000 238.880000 ;
      RECT 148.620000 237.800000 191.820000 238.880000 ;
      RECT 103.620000 237.800000 146.820000 238.880000 ;
      RECT 58.620000 237.800000 101.820000 238.880000 ;
      RECT 13.620000 237.800000 56.820000 238.880000 ;
      RECT 7.060000 237.800000 11.820000 238.880000 ;
      RECT 0.000000 237.800000 5.260000 238.880000 ;
      RECT 0.000000 237.440000 550.160000 237.800000 ;
      RECT 0.000000 236.460000 548.960000 237.440000 ;
      RECT 0.000000 236.160000 550.160000 236.460000 ;
      RECT 547.100000 235.080000 550.160000 236.160000 ;
      RECT 506.620000 235.080000 545.300000 236.160000 ;
      RECT 461.620000 235.080000 504.820000 236.160000 ;
      RECT 416.620000 235.080000 459.820000 236.160000 ;
      RECT 371.620000 235.080000 414.820000 236.160000 ;
      RECT 326.620000 235.080000 369.820000 236.160000 ;
      RECT 281.620000 235.080000 324.820000 236.160000 ;
      RECT 236.620000 235.080000 279.820000 236.160000 ;
      RECT 191.620000 235.080000 234.820000 236.160000 ;
      RECT 146.620000 235.080000 189.820000 236.160000 ;
      RECT 101.620000 235.080000 144.820000 236.160000 ;
      RECT 56.620000 235.080000 99.820000 236.160000 ;
      RECT 11.620000 235.080000 54.820000 236.160000 ;
      RECT 4.860000 235.080000 9.655000 236.160000 ;
      RECT 0.000000 235.080000 3.060000 236.160000 ;
      RECT 0.000000 233.780000 550.160000 235.080000 ;
      RECT 0.000000 233.440000 548.960000 233.780000 ;
      RECT 544.900000 232.800000 548.960000 233.440000 ;
      RECT 544.900000 232.360000 550.160000 232.800000 ;
      RECT 508.620000 232.360000 543.100000 233.440000 ;
      RECT 463.620000 232.360000 506.820000 233.440000 ;
      RECT 418.620000 232.360000 461.820000 233.440000 ;
      RECT 373.620000 232.360000 416.820000 233.440000 ;
      RECT 328.620000 232.360000 371.820000 233.440000 ;
      RECT 283.620000 232.360000 326.820000 233.440000 ;
      RECT 238.620000 232.360000 281.820000 233.440000 ;
      RECT 193.620000 232.360000 236.820000 233.440000 ;
      RECT 148.620000 232.360000 191.820000 233.440000 ;
      RECT 103.620000 232.360000 146.820000 233.440000 ;
      RECT 58.620000 232.360000 101.820000 233.440000 ;
      RECT 13.620000 232.360000 56.820000 233.440000 ;
      RECT 7.060000 232.360000 11.820000 233.440000 ;
      RECT 0.000000 232.360000 5.260000 233.440000 ;
      RECT 0.000000 230.730000 550.160000 232.360000 ;
      RECT 0.000000 230.720000 548.960000 230.730000 ;
      RECT 547.100000 229.750000 548.960000 230.720000 ;
      RECT 547.100000 229.640000 550.160000 229.750000 ;
      RECT 506.620000 229.640000 545.300000 230.720000 ;
      RECT 461.620000 229.640000 504.820000 230.720000 ;
      RECT 416.620000 229.640000 459.820000 230.720000 ;
      RECT 371.620000 229.640000 414.820000 230.720000 ;
      RECT 326.620000 229.640000 369.820000 230.720000 ;
      RECT 281.620000 229.640000 324.820000 230.720000 ;
      RECT 236.620000 229.640000 279.820000 230.720000 ;
      RECT 191.620000 229.640000 234.820000 230.720000 ;
      RECT 146.620000 229.640000 189.820000 230.720000 ;
      RECT 101.620000 229.640000 144.820000 230.720000 ;
      RECT 56.620000 229.640000 99.820000 230.720000 ;
      RECT 11.620000 229.640000 54.820000 230.720000 ;
      RECT 4.860000 229.640000 9.655000 230.720000 ;
      RECT 0.000000 229.640000 3.060000 230.720000 ;
      RECT 0.000000 228.000000 550.160000 229.640000 ;
      RECT 544.900000 227.680000 550.160000 228.000000 ;
      RECT 544.900000 226.920000 548.960000 227.680000 ;
      RECT 508.620000 226.920000 543.100000 228.000000 ;
      RECT 463.620000 226.920000 506.820000 228.000000 ;
      RECT 418.620000 226.920000 461.820000 228.000000 ;
      RECT 373.620000 226.920000 416.820000 228.000000 ;
      RECT 328.620000 226.920000 371.820000 228.000000 ;
      RECT 283.620000 226.920000 326.820000 228.000000 ;
      RECT 238.620000 226.920000 281.820000 228.000000 ;
      RECT 193.620000 226.920000 236.820000 228.000000 ;
      RECT 148.620000 226.920000 191.820000 228.000000 ;
      RECT 103.620000 226.920000 146.820000 228.000000 ;
      RECT 58.620000 226.920000 101.820000 228.000000 ;
      RECT 13.620000 226.920000 56.820000 228.000000 ;
      RECT 7.060000 226.920000 11.820000 228.000000 ;
      RECT 0.000000 226.920000 5.260000 228.000000 ;
      RECT 0.000000 226.700000 548.960000 226.920000 ;
      RECT 0.000000 225.280000 550.160000 226.700000 ;
      RECT 547.100000 224.630000 550.160000 225.280000 ;
      RECT 547.100000 224.200000 548.960000 224.630000 ;
      RECT 506.620000 224.200000 545.300000 225.280000 ;
      RECT 461.620000 224.200000 504.820000 225.280000 ;
      RECT 416.620000 224.200000 459.820000 225.280000 ;
      RECT 371.620000 224.200000 414.820000 225.280000 ;
      RECT 326.620000 224.200000 369.820000 225.280000 ;
      RECT 281.620000 224.200000 324.820000 225.280000 ;
      RECT 236.620000 224.200000 279.820000 225.280000 ;
      RECT 191.620000 224.200000 234.820000 225.280000 ;
      RECT 146.620000 224.200000 189.820000 225.280000 ;
      RECT 101.620000 224.200000 144.820000 225.280000 ;
      RECT 56.620000 224.200000 99.820000 225.280000 ;
      RECT 11.620000 224.200000 54.820000 225.280000 ;
      RECT 4.860000 224.200000 9.655000 225.280000 ;
      RECT 0.000000 224.200000 3.060000 225.280000 ;
      RECT 0.000000 223.650000 548.960000 224.200000 ;
      RECT 0.000000 222.560000 550.160000 223.650000 ;
      RECT 544.900000 221.580000 550.160000 222.560000 ;
      RECT 544.900000 221.480000 548.960000 221.580000 ;
      RECT 508.620000 221.480000 543.100000 222.560000 ;
      RECT 463.620000 221.480000 506.820000 222.560000 ;
      RECT 418.620000 221.480000 461.820000 222.560000 ;
      RECT 373.620000 221.480000 416.820000 222.560000 ;
      RECT 328.620000 221.480000 371.820000 222.560000 ;
      RECT 283.620000 221.480000 326.820000 222.560000 ;
      RECT 238.620000 221.480000 281.820000 222.560000 ;
      RECT 193.620000 221.480000 236.820000 222.560000 ;
      RECT 148.620000 221.480000 191.820000 222.560000 ;
      RECT 103.620000 221.480000 146.820000 222.560000 ;
      RECT 58.620000 221.480000 101.820000 222.560000 ;
      RECT 13.620000 221.480000 56.820000 222.560000 ;
      RECT 7.060000 221.480000 11.820000 222.560000 ;
      RECT 0.000000 221.480000 5.260000 222.560000 ;
      RECT 0.000000 220.600000 548.960000 221.480000 ;
      RECT 0.000000 219.840000 550.160000 220.600000 ;
      RECT 547.100000 218.760000 550.160000 219.840000 ;
      RECT 506.620000 218.760000 545.300000 219.840000 ;
      RECT 461.620000 218.760000 504.820000 219.840000 ;
      RECT 416.620000 218.760000 459.820000 219.840000 ;
      RECT 371.620000 218.760000 414.820000 219.840000 ;
      RECT 326.620000 218.760000 369.820000 219.840000 ;
      RECT 281.620000 218.760000 324.820000 219.840000 ;
      RECT 236.620000 218.760000 279.820000 219.840000 ;
      RECT 191.620000 218.760000 234.820000 219.840000 ;
      RECT 146.620000 218.760000 189.820000 219.840000 ;
      RECT 101.620000 218.760000 144.820000 219.840000 ;
      RECT 56.620000 218.760000 99.820000 219.840000 ;
      RECT 11.620000 218.760000 54.820000 219.840000 ;
      RECT 4.860000 218.760000 9.655000 219.840000 ;
      RECT 0.000000 218.760000 3.060000 219.840000 ;
      RECT 0.000000 218.530000 550.160000 218.760000 ;
      RECT 0.000000 217.550000 548.960000 218.530000 ;
      RECT 0.000000 217.120000 550.160000 217.550000 ;
      RECT 544.900000 216.040000 550.160000 217.120000 ;
      RECT 508.620000 216.040000 543.100000 217.120000 ;
      RECT 463.620000 216.040000 506.820000 217.120000 ;
      RECT 418.620000 216.040000 461.820000 217.120000 ;
      RECT 373.620000 216.040000 416.820000 217.120000 ;
      RECT 328.620000 216.040000 371.820000 217.120000 ;
      RECT 283.620000 216.040000 326.820000 217.120000 ;
      RECT 238.620000 216.040000 281.820000 217.120000 ;
      RECT 193.620000 216.040000 236.820000 217.120000 ;
      RECT 148.620000 216.040000 191.820000 217.120000 ;
      RECT 103.620000 216.040000 146.820000 217.120000 ;
      RECT 58.620000 216.040000 101.820000 217.120000 ;
      RECT 13.620000 216.040000 56.820000 217.120000 ;
      RECT 7.060000 216.040000 11.820000 217.120000 ;
      RECT 0.000000 216.040000 5.260000 217.120000 ;
      RECT 0.000000 214.870000 550.160000 216.040000 ;
      RECT 0.000000 214.400000 548.960000 214.870000 ;
      RECT 547.100000 213.890000 548.960000 214.400000 ;
      RECT 547.100000 213.320000 550.160000 213.890000 ;
      RECT 506.620000 213.320000 545.300000 214.400000 ;
      RECT 461.620000 213.320000 504.820000 214.400000 ;
      RECT 416.620000 213.320000 459.820000 214.400000 ;
      RECT 371.620000 213.320000 414.820000 214.400000 ;
      RECT 326.620000 213.320000 369.820000 214.400000 ;
      RECT 281.620000 213.320000 324.820000 214.400000 ;
      RECT 236.620000 213.320000 279.820000 214.400000 ;
      RECT 191.620000 213.320000 234.820000 214.400000 ;
      RECT 146.620000 213.320000 189.820000 214.400000 ;
      RECT 101.620000 213.320000 144.820000 214.400000 ;
      RECT 56.620000 213.320000 99.820000 214.400000 ;
      RECT 11.620000 213.320000 54.820000 214.400000 ;
      RECT 4.860000 213.320000 9.655000 214.400000 ;
      RECT 0.000000 213.320000 3.060000 214.400000 ;
      RECT 0.000000 211.820000 550.160000 213.320000 ;
      RECT 0.000000 211.680000 548.960000 211.820000 ;
      RECT 544.900000 210.840000 548.960000 211.680000 ;
      RECT 544.900000 210.600000 550.160000 210.840000 ;
      RECT 508.620000 210.600000 543.100000 211.680000 ;
      RECT 463.620000 210.600000 506.820000 211.680000 ;
      RECT 418.620000 210.600000 461.820000 211.680000 ;
      RECT 373.620000 210.600000 416.820000 211.680000 ;
      RECT 328.620000 210.600000 371.820000 211.680000 ;
      RECT 283.620000 210.600000 326.820000 211.680000 ;
      RECT 238.620000 210.600000 281.820000 211.680000 ;
      RECT 193.620000 210.600000 236.820000 211.680000 ;
      RECT 148.620000 210.600000 191.820000 211.680000 ;
      RECT 103.620000 210.600000 146.820000 211.680000 ;
      RECT 58.620000 210.600000 101.820000 211.680000 ;
      RECT 13.620000 210.600000 56.820000 211.680000 ;
      RECT 7.060000 210.600000 11.820000 211.680000 ;
      RECT 0.000000 210.600000 5.260000 211.680000 ;
      RECT 0.000000 208.960000 550.160000 210.600000 ;
      RECT 547.100000 208.770000 550.160000 208.960000 ;
      RECT 547.100000 207.880000 548.960000 208.770000 ;
      RECT 506.620000 207.880000 545.300000 208.960000 ;
      RECT 461.620000 207.880000 504.820000 208.960000 ;
      RECT 416.620000 207.880000 459.820000 208.960000 ;
      RECT 371.620000 207.880000 414.820000 208.960000 ;
      RECT 326.620000 207.880000 369.820000 208.960000 ;
      RECT 281.620000 207.880000 324.820000 208.960000 ;
      RECT 236.620000 207.880000 279.820000 208.960000 ;
      RECT 191.620000 207.880000 234.820000 208.960000 ;
      RECT 146.620000 207.880000 189.820000 208.960000 ;
      RECT 101.620000 207.880000 144.820000 208.960000 ;
      RECT 56.620000 207.880000 99.820000 208.960000 ;
      RECT 11.620000 207.880000 54.820000 208.960000 ;
      RECT 4.860000 207.880000 9.655000 208.960000 ;
      RECT 0.000000 207.880000 3.060000 208.960000 ;
      RECT 0.000000 207.790000 548.960000 207.880000 ;
      RECT 0.000000 206.240000 550.160000 207.790000 ;
      RECT 544.900000 205.720000 550.160000 206.240000 ;
      RECT 544.900000 205.160000 548.960000 205.720000 ;
      RECT 508.620000 205.160000 543.100000 206.240000 ;
      RECT 463.620000 205.160000 506.820000 206.240000 ;
      RECT 418.620000 205.160000 461.820000 206.240000 ;
      RECT 373.620000 205.160000 416.820000 206.240000 ;
      RECT 328.620000 205.160000 371.820000 206.240000 ;
      RECT 283.620000 205.160000 326.820000 206.240000 ;
      RECT 238.620000 205.160000 281.820000 206.240000 ;
      RECT 193.620000 205.160000 236.820000 206.240000 ;
      RECT 148.620000 205.160000 191.820000 206.240000 ;
      RECT 103.620000 205.160000 146.820000 206.240000 ;
      RECT 58.620000 205.160000 101.820000 206.240000 ;
      RECT 13.620000 205.160000 56.820000 206.240000 ;
      RECT 7.060000 205.160000 11.820000 206.240000 ;
      RECT 0.000000 205.160000 5.260000 206.240000 ;
      RECT 0.000000 204.740000 548.960000 205.160000 ;
      RECT 0.000000 203.520000 550.160000 204.740000 ;
      RECT 547.100000 202.670000 550.160000 203.520000 ;
      RECT 547.100000 202.440000 548.960000 202.670000 ;
      RECT 506.620000 202.440000 545.300000 203.520000 ;
      RECT 461.620000 202.440000 504.820000 203.520000 ;
      RECT 416.620000 202.440000 459.820000 203.520000 ;
      RECT 371.620000 202.440000 414.820000 203.520000 ;
      RECT 326.620000 202.440000 369.820000 203.520000 ;
      RECT 281.620000 202.440000 324.820000 203.520000 ;
      RECT 236.620000 202.440000 279.820000 203.520000 ;
      RECT 191.620000 202.440000 234.820000 203.520000 ;
      RECT 146.620000 202.440000 189.820000 203.520000 ;
      RECT 101.620000 202.440000 144.820000 203.520000 ;
      RECT 56.620000 202.440000 99.820000 203.520000 ;
      RECT 11.620000 202.440000 54.820000 203.520000 ;
      RECT 4.860000 202.440000 9.655000 203.520000 ;
      RECT 0.000000 202.440000 3.060000 203.520000 ;
      RECT 0.000000 201.690000 548.960000 202.440000 ;
      RECT 0.000000 200.800000 550.160000 201.690000 ;
      RECT 544.900000 199.720000 550.160000 200.800000 ;
      RECT 508.620000 199.720000 543.100000 200.800000 ;
      RECT 463.620000 199.720000 506.820000 200.800000 ;
      RECT 418.620000 199.720000 461.820000 200.800000 ;
      RECT 373.620000 199.720000 416.820000 200.800000 ;
      RECT 328.620000 199.720000 371.820000 200.800000 ;
      RECT 283.620000 199.720000 326.820000 200.800000 ;
      RECT 238.620000 199.720000 281.820000 200.800000 ;
      RECT 193.620000 199.720000 236.820000 200.800000 ;
      RECT 148.620000 199.720000 191.820000 200.800000 ;
      RECT 103.620000 199.720000 146.820000 200.800000 ;
      RECT 58.620000 199.720000 101.820000 200.800000 ;
      RECT 13.620000 199.720000 56.820000 200.800000 ;
      RECT 7.060000 199.720000 11.820000 200.800000 ;
      RECT 0.000000 199.720000 5.260000 200.800000 ;
      RECT 0.000000 199.620000 550.160000 199.720000 ;
      RECT 0.000000 198.640000 548.960000 199.620000 ;
      RECT 0.000000 198.080000 550.160000 198.640000 ;
      RECT 547.100000 197.000000 550.160000 198.080000 ;
      RECT 506.620000 197.000000 545.300000 198.080000 ;
      RECT 461.620000 197.000000 504.820000 198.080000 ;
      RECT 416.620000 197.000000 459.820000 198.080000 ;
      RECT 371.620000 197.000000 414.820000 198.080000 ;
      RECT 326.620000 197.000000 369.820000 198.080000 ;
      RECT 281.620000 197.000000 324.820000 198.080000 ;
      RECT 236.620000 197.000000 279.820000 198.080000 ;
      RECT 191.620000 197.000000 234.820000 198.080000 ;
      RECT 146.620000 197.000000 189.820000 198.080000 ;
      RECT 101.620000 197.000000 144.820000 198.080000 ;
      RECT 56.620000 197.000000 99.820000 198.080000 ;
      RECT 11.620000 197.000000 54.820000 198.080000 ;
      RECT 4.860000 197.000000 9.655000 198.080000 ;
      RECT 0.000000 197.000000 3.060000 198.080000 ;
      RECT 0.000000 195.960000 550.160000 197.000000 ;
      RECT 0.000000 195.360000 548.960000 195.960000 ;
      RECT 544.900000 194.980000 548.960000 195.360000 ;
      RECT 544.900000 194.280000 550.160000 194.980000 ;
      RECT 508.620000 194.280000 543.100000 195.360000 ;
      RECT 463.620000 194.280000 506.820000 195.360000 ;
      RECT 418.620000 194.280000 461.820000 195.360000 ;
      RECT 373.620000 194.280000 416.820000 195.360000 ;
      RECT 328.620000 194.280000 371.820000 195.360000 ;
      RECT 283.620000 194.280000 326.820000 195.360000 ;
      RECT 238.620000 194.280000 281.820000 195.360000 ;
      RECT 193.620000 194.280000 236.820000 195.360000 ;
      RECT 148.620000 194.280000 191.820000 195.360000 ;
      RECT 103.620000 194.280000 146.820000 195.360000 ;
      RECT 58.620000 194.280000 101.820000 195.360000 ;
      RECT 13.620000 194.280000 56.820000 195.360000 ;
      RECT 7.060000 194.280000 11.820000 195.360000 ;
      RECT 0.000000 194.280000 5.260000 195.360000 ;
      RECT 0.000000 192.910000 550.160000 194.280000 ;
      RECT 0.000000 192.640000 548.960000 192.910000 ;
      RECT 547.100000 191.930000 548.960000 192.640000 ;
      RECT 547.100000 191.560000 550.160000 191.930000 ;
      RECT 506.620000 191.560000 545.300000 192.640000 ;
      RECT 461.620000 191.560000 504.820000 192.640000 ;
      RECT 416.620000 191.560000 459.820000 192.640000 ;
      RECT 371.620000 191.560000 414.820000 192.640000 ;
      RECT 326.620000 191.560000 369.820000 192.640000 ;
      RECT 281.620000 191.560000 324.820000 192.640000 ;
      RECT 236.620000 191.560000 279.820000 192.640000 ;
      RECT 191.620000 191.560000 234.820000 192.640000 ;
      RECT 146.620000 191.560000 189.820000 192.640000 ;
      RECT 101.620000 191.560000 144.820000 192.640000 ;
      RECT 56.620000 191.560000 99.820000 192.640000 ;
      RECT 11.620000 191.560000 54.820000 192.640000 ;
      RECT 4.860000 191.560000 9.655000 192.640000 ;
      RECT 0.000000 191.560000 3.060000 192.640000 ;
      RECT 0.000000 189.920000 550.160000 191.560000 ;
      RECT 544.900000 189.860000 550.160000 189.920000 ;
      RECT 544.900000 188.880000 548.960000 189.860000 ;
      RECT 544.900000 188.840000 550.160000 188.880000 ;
      RECT 508.620000 188.840000 543.100000 189.920000 ;
      RECT 463.620000 188.840000 506.820000 189.920000 ;
      RECT 418.620000 188.840000 461.820000 189.920000 ;
      RECT 373.620000 188.840000 416.820000 189.920000 ;
      RECT 328.620000 188.840000 371.820000 189.920000 ;
      RECT 283.620000 188.840000 326.820000 189.920000 ;
      RECT 238.620000 188.840000 281.820000 189.920000 ;
      RECT 193.620000 188.840000 236.820000 189.920000 ;
      RECT 148.620000 188.840000 191.820000 189.920000 ;
      RECT 103.620000 188.840000 146.820000 189.920000 ;
      RECT 58.620000 188.840000 101.820000 189.920000 ;
      RECT 13.620000 188.840000 56.820000 189.920000 ;
      RECT 7.060000 188.840000 11.820000 189.920000 ;
      RECT 0.000000 188.840000 5.260000 189.920000 ;
      RECT 0.000000 187.200000 550.160000 188.840000 ;
      RECT 547.100000 186.810000 550.160000 187.200000 ;
      RECT 547.100000 186.120000 548.960000 186.810000 ;
      RECT 506.620000 186.120000 545.300000 187.200000 ;
      RECT 461.620000 186.120000 504.820000 187.200000 ;
      RECT 416.620000 186.120000 459.820000 187.200000 ;
      RECT 371.620000 186.120000 414.820000 187.200000 ;
      RECT 326.620000 186.120000 369.820000 187.200000 ;
      RECT 281.620000 186.120000 324.820000 187.200000 ;
      RECT 236.620000 186.120000 279.820000 187.200000 ;
      RECT 191.620000 186.120000 234.820000 187.200000 ;
      RECT 146.620000 186.120000 189.820000 187.200000 ;
      RECT 101.620000 186.120000 144.820000 187.200000 ;
      RECT 56.620000 186.120000 99.820000 187.200000 ;
      RECT 11.620000 186.120000 54.820000 187.200000 ;
      RECT 4.860000 186.120000 9.655000 187.200000 ;
      RECT 0.000000 186.120000 3.060000 187.200000 ;
      RECT 0.000000 185.830000 548.960000 186.120000 ;
      RECT 0.000000 184.480000 550.160000 185.830000 ;
      RECT 544.900000 183.760000 550.160000 184.480000 ;
      RECT 544.900000 183.400000 548.960000 183.760000 ;
      RECT 508.620000 183.400000 543.100000 184.480000 ;
      RECT 463.620000 183.400000 506.820000 184.480000 ;
      RECT 418.620000 183.400000 461.820000 184.480000 ;
      RECT 373.620000 183.400000 416.820000 184.480000 ;
      RECT 328.620000 183.400000 371.820000 184.480000 ;
      RECT 283.620000 183.400000 326.820000 184.480000 ;
      RECT 238.620000 183.400000 281.820000 184.480000 ;
      RECT 193.620000 183.400000 236.820000 184.480000 ;
      RECT 148.620000 183.400000 191.820000 184.480000 ;
      RECT 103.620000 183.400000 146.820000 184.480000 ;
      RECT 58.620000 183.400000 101.820000 184.480000 ;
      RECT 13.620000 183.400000 56.820000 184.480000 ;
      RECT 7.060000 183.400000 11.820000 184.480000 ;
      RECT 0.000000 183.400000 5.260000 184.480000 ;
      RECT 0.000000 182.780000 548.960000 183.400000 ;
      RECT 0.000000 181.760000 550.160000 182.780000 ;
      RECT 547.100000 180.680000 550.160000 181.760000 ;
      RECT 506.620000 180.680000 545.300000 181.760000 ;
      RECT 461.620000 180.680000 504.820000 181.760000 ;
      RECT 416.620000 180.680000 459.820000 181.760000 ;
      RECT 371.620000 180.680000 414.820000 181.760000 ;
      RECT 326.620000 180.680000 369.820000 181.760000 ;
      RECT 281.620000 180.680000 324.820000 181.760000 ;
      RECT 236.620000 180.680000 279.820000 181.760000 ;
      RECT 191.620000 180.680000 234.820000 181.760000 ;
      RECT 146.620000 180.680000 189.820000 181.760000 ;
      RECT 101.620000 180.680000 144.820000 181.760000 ;
      RECT 56.620000 180.680000 99.820000 181.760000 ;
      RECT 11.620000 180.680000 54.820000 181.760000 ;
      RECT 4.860000 180.680000 9.655000 181.760000 ;
      RECT 0.000000 180.680000 3.060000 181.760000 ;
      RECT 0.000000 180.100000 550.160000 180.680000 ;
      RECT 0.000000 179.120000 548.960000 180.100000 ;
      RECT 0.000000 179.040000 550.160000 179.120000 ;
      RECT 544.900000 177.960000 550.160000 179.040000 ;
      RECT 508.620000 177.960000 543.100000 179.040000 ;
      RECT 463.620000 177.960000 506.820000 179.040000 ;
      RECT 418.620000 177.960000 461.820000 179.040000 ;
      RECT 373.620000 177.960000 416.820000 179.040000 ;
      RECT 328.620000 177.960000 371.820000 179.040000 ;
      RECT 283.620000 177.960000 326.820000 179.040000 ;
      RECT 238.620000 177.960000 281.820000 179.040000 ;
      RECT 193.620000 177.960000 236.820000 179.040000 ;
      RECT 148.620000 177.960000 191.820000 179.040000 ;
      RECT 103.620000 177.960000 146.820000 179.040000 ;
      RECT 58.620000 177.960000 101.820000 179.040000 ;
      RECT 13.620000 177.960000 56.820000 179.040000 ;
      RECT 7.060000 177.960000 11.820000 179.040000 ;
      RECT 0.000000 177.960000 5.260000 179.040000 ;
      RECT 0.000000 177.050000 550.160000 177.960000 ;
      RECT 0.000000 176.320000 548.960000 177.050000 ;
      RECT 547.100000 176.070000 548.960000 176.320000 ;
      RECT 547.100000 175.240000 550.160000 176.070000 ;
      RECT 506.620000 175.240000 545.300000 176.320000 ;
      RECT 461.620000 175.240000 504.820000 176.320000 ;
      RECT 416.620000 175.240000 459.820000 176.320000 ;
      RECT 371.620000 175.240000 414.820000 176.320000 ;
      RECT 326.620000 175.240000 369.820000 176.320000 ;
      RECT 281.620000 175.240000 324.820000 176.320000 ;
      RECT 236.620000 175.240000 279.820000 176.320000 ;
      RECT 191.620000 175.240000 234.820000 176.320000 ;
      RECT 146.620000 175.240000 189.820000 176.320000 ;
      RECT 101.620000 175.240000 144.820000 176.320000 ;
      RECT 56.620000 175.240000 99.820000 176.320000 ;
      RECT 11.620000 175.240000 54.820000 176.320000 ;
      RECT 4.860000 175.240000 9.655000 176.320000 ;
      RECT 0.000000 175.240000 3.060000 176.320000 ;
      RECT 0.000000 174.000000 550.160000 175.240000 ;
      RECT 0.000000 173.600000 548.960000 174.000000 ;
      RECT 544.900000 173.020000 548.960000 173.600000 ;
      RECT 544.900000 172.520000 550.160000 173.020000 ;
      RECT 508.620000 172.520000 543.100000 173.600000 ;
      RECT 463.620000 172.520000 506.820000 173.600000 ;
      RECT 418.620000 172.520000 461.820000 173.600000 ;
      RECT 373.620000 172.520000 416.820000 173.600000 ;
      RECT 328.620000 172.520000 371.820000 173.600000 ;
      RECT 283.620000 172.520000 326.820000 173.600000 ;
      RECT 238.620000 172.520000 281.820000 173.600000 ;
      RECT 193.620000 172.520000 236.820000 173.600000 ;
      RECT 148.620000 172.520000 191.820000 173.600000 ;
      RECT 103.620000 172.520000 146.820000 173.600000 ;
      RECT 58.620000 172.520000 101.820000 173.600000 ;
      RECT 13.620000 172.520000 56.820000 173.600000 ;
      RECT 7.060000 172.520000 11.820000 173.600000 ;
      RECT 0.000000 172.520000 5.260000 173.600000 ;
      RECT 0.000000 170.950000 550.160000 172.520000 ;
      RECT 0.000000 170.880000 548.960000 170.950000 ;
      RECT 547.100000 169.970000 548.960000 170.880000 ;
      RECT 547.100000 169.800000 550.160000 169.970000 ;
      RECT 506.620000 169.800000 545.300000 170.880000 ;
      RECT 461.620000 169.800000 504.820000 170.880000 ;
      RECT 416.620000 169.800000 459.820000 170.880000 ;
      RECT 371.620000 169.800000 414.820000 170.880000 ;
      RECT 326.620000 169.800000 369.820000 170.880000 ;
      RECT 281.620000 169.800000 324.820000 170.880000 ;
      RECT 236.620000 169.800000 279.820000 170.880000 ;
      RECT 191.620000 169.800000 234.820000 170.880000 ;
      RECT 146.620000 169.800000 189.820000 170.880000 ;
      RECT 101.620000 169.800000 144.820000 170.880000 ;
      RECT 56.620000 169.800000 99.820000 170.880000 ;
      RECT 11.620000 169.800000 54.820000 170.880000 ;
      RECT 4.860000 169.800000 9.655000 170.880000 ;
      RECT 0.000000 169.800000 3.060000 170.880000 ;
      RECT 0.000000 168.160000 550.160000 169.800000 ;
      RECT 544.900000 167.900000 550.160000 168.160000 ;
      RECT 544.900000 167.080000 548.960000 167.900000 ;
      RECT 508.620000 167.080000 543.100000 168.160000 ;
      RECT 463.620000 167.080000 506.820000 168.160000 ;
      RECT 418.620000 167.080000 461.820000 168.160000 ;
      RECT 373.620000 167.080000 416.820000 168.160000 ;
      RECT 328.620000 167.080000 371.820000 168.160000 ;
      RECT 283.620000 167.080000 326.820000 168.160000 ;
      RECT 238.620000 167.080000 281.820000 168.160000 ;
      RECT 193.620000 167.080000 236.820000 168.160000 ;
      RECT 148.620000 167.080000 191.820000 168.160000 ;
      RECT 103.620000 167.080000 146.820000 168.160000 ;
      RECT 58.620000 167.080000 101.820000 168.160000 ;
      RECT 13.620000 167.080000 56.820000 168.160000 ;
      RECT 7.060000 167.080000 11.820000 168.160000 ;
      RECT 0.000000 167.080000 5.260000 168.160000 ;
      RECT 0.000000 166.920000 548.960000 167.080000 ;
      RECT 0.000000 165.440000 550.160000 166.920000 ;
      RECT 547.100000 164.850000 550.160000 165.440000 ;
      RECT 547.100000 164.360000 548.960000 164.850000 ;
      RECT 506.620000 164.360000 545.300000 165.440000 ;
      RECT 461.620000 164.360000 504.820000 165.440000 ;
      RECT 416.620000 164.360000 459.820000 165.440000 ;
      RECT 371.620000 164.360000 414.820000 165.440000 ;
      RECT 326.620000 164.360000 369.820000 165.440000 ;
      RECT 281.620000 164.360000 324.820000 165.440000 ;
      RECT 236.620000 164.360000 279.820000 165.440000 ;
      RECT 191.620000 164.360000 234.820000 165.440000 ;
      RECT 146.620000 164.360000 189.820000 165.440000 ;
      RECT 101.620000 164.360000 144.820000 165.440000 ;
      RECT 56.620000 164.360000 99.820000 165.440000 ;
      RECT 11.620000 164.360000 54.820000 165.440000 ;
      RECT 4.860000 164.360000 9.655000 165.440000 ;
      RECT 0.000000 164.360000 3.060000 165.440000 ;
      RECT 0.000000 163.870000 548.960000 164.360000 ;
      RECT 0.000000 162.720000 550.160000 163.870000 ;
      RECT 544.900000 161.640000 550.160000 162.720000 ;
      RECT 508.620000 161.640000 543.100000 162.720000 ;
      RECT 463.620000 161.640000 506.820000 162.720000 ;
      RECT 418.620000 161.640000 461.820000 162.720000 ;
      RECT 373.620000 161.640000 416.820000 162.720000 ;
      RECT 328.620000 161.640000 371.820000 162.720000 ;
      RECT 283.620000 161.640000 326.820000 162.720000 ;
      RECT 238.620000 161.640000 281.820000 162.720000 ;
      RECT 193.620000 161.640000 236.820000 162.720000 ;
      RECT 148.620000 161.640000 191.820000 162.720000 ;
      RECT 103.620000 161.640000 146.820000 162.720000 ;
      RECT 58.620000 161.640000 101.820000 162.720000 ;
      RECT 13.620000 161.640000 56.820000 162.720000 ;
      RECT 7.060000 161.640000 11.820000 162.720000 ;
      RECT 0.000000 161.640000 5.260000 162.720000 ;
      RECT 0.000000 161.190000 550.160000 161.640000 ;
      RECT 0.000000 160.210000 548.960000 161.190000 ;
      RECT 0.000000 160.000000 550.160000 160.210000 ;
      RECT 547.100000 158.920000 550.160000 160.000000 ;
      RECT 506.620000 158.920000 545.300000 160.000000 ;
      RECT 461.620000 158.920000 504.820000 160.000000 ;
      RECT 416.620000 158.920000 459.820000 160.000000 ;
      RECT 371.620000 158.920000 414.820000 160.000000 ;
      RECT 326.620000 158.920000 369.820000 160.000000 ;
      RECT 281.620000 158.920000 324.820000 160.000000 ;
      RECT 236.620000 158.920000 279.820000 160.000000 ;
      RECT 191.620000 158.920000 234.820000 160.000000 ;
      RECT 146.620000 158.920000 189.820000 160.000000 ;
      RECT 101.620000 158.920000 144.820000 160.000000 ;
      RECT 56.620000 158.920000 99.820000 160.000000 ;
      RECT 11.620000 158.920000 54.820000 160.000000 ;
      RECT 4.860000 158.920000 9.655000 160.000000 ;
      RECT 0.000000 158.920000 3.060000 160.000000 ;
      RECT 0.000000 158.140000 550.160000 158.920000 ;
      RECT 0.000000 157.280000 548.960000 158.140000 ;
      RECT 544.900000 157.160000 548.960000 157.280000 ;
      RECT 544.900000 156.200000 550.160000 157.160000 ;
      RECT 508.620000 156.200000 543.100000 157.280000 ;
      RECT 463.620000 156.200000 506.820000 157.280000 ;
      RECT 418.620000 156.200000 461.820000 157.280000 ;
      RECT 373.620000 156.200000 416.820000 157.280000 ;
      RECT 328.620000 156.200000 371.820000 157.280000 ;
      RECT 283.620000 156.200000 326.820000 157.280000 ;
      RECT 238.620000 156.200000 281.820000 157.280000 ;
      RECT 193.620000 156.200000 236.820000 157.280000 ;
      RECT 148.620000 156.200000 191.820000 157.280000 ;
      RECT 103.620000 156.200000 146.820000 157.280000 ;
      RECT 58.620000 156.200000 101.820000 157.280000 ;
      RECT 13.620000 156.200000 56.820000 157.280000 ;
      RECT 7.060000 156.200000 11.820000 157.280000 ;
      RECT 0.000000 156.200000 5.260000 157.280000 ;
      RECT 0.000000 155.090000 550.160000 156.200000 ;
      RECT 0.000000 154.560000 548.960000 155.090000 ;
      RECT 547.100000 154.110000 548.960000 154.560000 ;
      RECT 547.100000 153.480000 550.160000 154.110000 ;
      RECT 506.620000 153.480000 545.300000 154.560000 ;
      RECT 461.620000 153.480000 504.820000 154.560000 ;
      RECT 416.620000 153.480000 459.820000 154.560000 ;
      RECT 371.620000 153.480000 414.820000 154.560000 ;
      RECT 326.620000 153.480000 369.820000 154.560000 ;
      RECT 281.620000 153.480000 324.820000 154.560000 ;
      RECT 236.620000 153.480000 279.820000 154.560000 ;
      RECT 191.620000 153.480000 234.820000 154.560000 ;
      RECT 146.620000 153.480000 189.820000 154.560000 ;
      RECT 101.620000 153.480000 144.820000 154.560000 ;
      RECT 56.620000 153.480000 99.820000 154.560000 ;
      RECT 11.620000 153.480000 54.820000 154.560000 ;
      RECT 4.860000 153.480000 9.655000 154.560000 ;
      RECT 0.000000 153.480000 3.060000 154.560000 ;
      RECT 0.000000 152.040000 550.160000 153.480000 ;
      RECT 0.000000 151.840000 548.960000 152.040000 ;
      RECT 544.900000 151.060000 548.960000 151.840000 ;
      RECT 544.900000 150.760000 550.160000 151.060000 ;
      RECT 508.620000 150.760000 543.100000 151.840000 ;
      RECT 463.620000 150.760000 506.820000 151.840000 ;
      RECT 418.620000 150.760000 461.820000 151.840000 ;
      RECT 373.620000 150.760000 416.820000 151.840000 ;
      RECT 328.620000 150.760000 371.820000 151.840000 ;
      RECT 283.620000 150.760000 326.820000 151.840000 ;
      RECT 238.620000 150.760000 281.820000 151.840000 ;
      RECT 193.620000 150.760000 236.820000 151.840000 ;
      RECT 148.620000 150.760000 191.820000 151.840000 ;
      RECT 103.620000 150.760000 146.820000 151.840000 ;
      RECT 58.620000 150.760000 101.820000 151.840000 ;
      RECT 13.620000 150.760000 56.820000 151.840000 ;
      RECT 7.060000 150.760000 11.820000 151.840000 ;
      RECT 0.000000 150.760000 5.260000 151.840000 ;
      RECT 0.000000 149.120000 550.160000 150.760000 ;
      RECT 547.100000 148.990000 550.160000 149.120000 ;
      RECT 547.100000 148.040000 548.960000 148.990000 ;
      RECT 506.620000 148.040000 545.300000 149.120000 ;
      RECT 461.620000 148.040000 504.820000 149.120000 ;
      RECT 416.620000 148.040000 459.820000 149.120000 ;
      RECT 371.620000 148.040000 414.820000 149.120000 ;
      RECT 326.620000 148.040000 369.820000 149.120000 ;
      RECT 281.620000 148.040000 324.820000 149.120000 ;
      RECT 236.620000 148.040000 279.820000 149.120000 ;
      RECT 191.620000 148.040000 234.820000 149.120000 ;
      RECT 146.620000 148.040000 189.820000 149.120000 ;
      RECT 101.620000 148.040000 144.820000 149.120000 ;
      RECT 56.620000 148.040000 99.820000 149.120000 ;
      RECT 11.620000 148.040000 54.820000 149.120000 ;
      RECT 4.860000 148.040000 9.655000 149.120000 ;
      RECT 0.000000 148.040000 3.060000 149.120000 ;
      RECT 0.000000 148.010000 548.960000 148.040000 ;
      RECT 0.000000 146.400000 550.160000 148.010000 ;
      RECT 544.900000 145.940000 550.160000 146.400000 ;
      RECT 544.900000 145.320000 548.960000 145.940000 ;
      RECT 508.620000 145.320000 543.100000 146.400000 ;
      RECT 463.620000 145.320000 506.820000 146.400000 ;
      RECT 418.620000 145.320000 461.820000 146.400000 ;
      RECT 373.620000 145.320000 416.820000 146.400000 ;
      RECT 328.620000 145.320000 371.820000 146.400000 ;
      RECT 283.620000 145.320000 326.820000 146.400000 ;
      RECT 238.620000 145.320000 281.820000 146.400000 ;
      RECT 193.620000 145.320000 236.820000 146.400000 ;
      RECT 148.620000 145.320000 191.820000 146.400000 ;
      RECT 103.620000 145.320000 146.820000 146.400000 ;
      RECT 58.620000 145.320000 101.820000 146.400000 ;
      RECT 13.620000 145.320000 56.820000 146.400000 ;
      RECT 7.060000 145.320000 11.820000 146.400000 ;
      RECT 0.000000 145.320000 5.260000 146.400000 ;
      RECT 0.000000 144.960000 548.960000 145.320000 ;
      RECT 0.000000 143.680000 550.160000 144.960000 ;
      RECT 547.100000 142.600000 550.160000 143.680000 ;
      RECT 506.620000 142.600000 545.300000 143.680000 ;
      RECT 461.620000 142.600000 504.820000 143.680000 ;
      RECT 416.620000 142.600000 459.820000 143.680000 ;
      RECT 371.620000 142.600000 414.820000 143.680000 ;
      RECT 326.620000 142.600000 369.820000 143.680000 ;
      RECT 281.620000 142.600000 324.820000 143.680000 ;
      RECT 236.620000 142.600000 279.820000 143.680000 ;
      RECT 191.620000 142.600000 234.820000 143.680000 ;
      RECT 146.620000 142.600000 189.820000 143.680000 ;
      RECT 101.620000 142.600000 144.820000 143.680000 ;
      RECT 56.620000 142.600000 99.820000 143.680000 ;
      RECT 11.620000 142.600000 54.820000 143.680000 ;
      RECT 4.860000 142.600000 9.655000 143.680000 ;
      RECT 0.000000 142.600000 3.060000 143.680000 ;
      RECT 0.000000 142.280000 550.160000 142.600000 ;
      RECT 0.000000 141.300000 548.960000 142.280000 ;
      RECT 0.000000 140.960000 550.160000 141.300000 ;
      RECT 544.900000 139.880000 550.160000 140.960000 ;
      RECT 508.620000 139.880000 543.100000 140.960000 ;
      RECT 463.620000 139.880000 506.820000 140.960000 ;
      RECT 418.620000 139.880000 461.820000 140.960000 ;
      RECT 373.620000 139.880000 416.820000 140.960000 ;
      RECT 328.620000 139.880000 371.820000 140.960000 ;
      RECT 283.620000 139.880000 326.820000 140.960000 ;
      RECT 238.620000 139.880000 281.820000 140.960000 ;
      RECT 193.620000 139.880000 236.820000 140.960000 ;
      RECT 148.620000 139.880000 191.820000 140.960000 ;
      RECT 103.620000 139.880000 146.820000 140.960000 ;
      RECT 58.620000 139.880000 101.820000 140.960000 ;
      RECT 13.620000 139.880000 56.820000 140.960000 ;
      RECT 7.060000 139.880000 11.820000 140.960000 ;
      RECT 0.000000 139.880000 5.260000 140.960000 ;
      RECT 0.000000 139.230000 550.160000 139.880000 ;
      RECT 0.000000 138.250000 548.960000 139.230000 ;
      RECT 0.000000 138.240000 550.160000 138.250000 ;
      RECT 547.100000 137.160000 550.160000 138.240000 ;
      RECT 506.620000 137.160000 545.300000 138.240000 ;
      RECT 461.620000 137.160000 504.820000 138.240000 ;
      RECT 416.620000 137.160000 459.820000 138.240000 ;
      RECT 371.620000 137.160000 414.820000 138.240000 ;
      RECT 326.620000 137.160000 369.820000 138.240000 ;
      RECT 281.620000 137.160000 324.820000 138.240000 ;
      RECT 236.620000 137.160000 279.820000 138.240000 ;
      RECT 191.620000 137.160000 234.820000 138.240000 ;
      RECT 146.620000 137.160000 189.820000 138.240000 ;
      RECT 101.620000 137.160000 144.820000 138.240000 ;
      RECT 56.620000 137.160000 99.820000 138.240000 ;
      RECT 11.620000 137.160000 54.820000 138.240000 ;
      RECT 4.860000 137.160000 9.655000 138.240000 ;
      RECT 0.000000 137.160000 3.060000 138.240000 ;
      RECT 0.000000 136.180000 550.160000 137.160000 ;
      RECT 0.000000 135.520000 548.960000 136.180000 ;
      RECT 544.900000 135.200000 548.960000 135.520000 ;
      RECT 544.900000 134.440000 550.160000 135.200000 ;
      RECT 508.620000 134.440000 543.100000 135.520000 ;
      RECT 463.620000 134.440000 506.820000 135.520000 ;
      RECT 418.620000 134.440000 461.820000 135.520000 ;
      RECT 373.620000 134.440000 416.820000 135.520000 ;
      RECT 328.620000 134.440000 371.820000 135.520000 ;
      RECT 283.620000 134.440000 326.820000 135.520000 ;
      RECT 238.620000 134.440000 281.820000 135.520000 ;
      RECT 193.620000 134.440000 236.820000 135.520000 ;
      RECT 148.620000 134.440000 191.820000 135.520000 ;
      RECT 103.620000 134.440000 146.820000 135.520000 ;
      RECT 58.620000 134.440000 101.820000 135.520000 ;
      RECT 13.620000 134.440000 56.820000 135.520000 ;
      RECT 7.060000 134.440000 11.820000 135.520000 ;
      RECT 0.000000 134.440000 5.260000 135.520000 ;
      RECT 0.000000 133.130000 550.160000 134.440000 ;
      RECT 0.000000 132.800000 548.960000 133.130000 ;
      RECT 547.100000 132.150000 548.960000 132.800000 ;
      RECT 547.100000 131.720000 550.160000 132.150000 ;
      RECT 506.620000 131.720000 545.300000 132.800000 ;
      RECT 461.620000 131.720000 504.820000 132.800000 ;
      RECT 416.620000 131.720000 459.820000 132.800000 ;
      RECT 371.620000 131.720000 414.820000 132.800000 ;
      RECT 326.620000 131.720000 369.820000 132.800000 ;
      RECT 281.620000 131.720000 324.820000 132.800000 ;
      RECT 236.620000 131.720000 279.820000 132.800000 ;
      RECT 191.620000 131.720000 234.820000 132.800000 ;
      RECT 146.620000 131.720000 189.820000 132.800000 ;
      RECT 101.620000 131.720000 144.820000 132.800000 ;
      RECT 56.620000 131.720000 99.820000 132.800000 ;
      RECT 11.620000 131.720000 54.820000 132.800000 ;
      RECT 4.860000 131.720000 9.655000 132.800000 ;
      RECT 0.000000 131.720000 3.060000 132.800000 ;
      RECT 0.000000 130.080000 550.160000 131.720000 ;
      RECT 544.900000 129.100000 548.960000 130.080000 ;
      RECT 544.900000 129.000000 550.160000 129.100000 ;
      RECT 508.620000 129.000000 543.100000 130.080000 ;
      RECT 463.620000 129.000000 506.820000 130.080000 ;
      RECT 418.620000 129.000000 461.820000 130.080000 ;
      RECT 373.620000 129.000000 416.820000 130.080000 ;
      RECT 328.620000 129.000000 371.820000 130.080000 ;
      RECT 283.620000 129.000000 326.820000 130.080000 ;
      RECT 238.620000 129.000000 281.820000 130.080000 ;
      RECT 193.620000 129.000000 236.820000 130.080000 ;
      RECT 148.620000 129.000000 191.820000 130.080000 ;
      RECT 103.620000 129.000000 146.820000 130.080000 ;
      RECT 58.620000 129.000000 101.820000 130.080000 ;
      RECT 13.620000 129.000000 56.820000 130.080000 ;
      RECT 7.060000 129.000000 11.820000 130.080000 ;
      RECT 0.000000 129.000000 5.260000 130.080000 ;
      RECT 0.000000 127.360000 550.160000 129.000000 ;
      RECT 547.100000 127.030000 550.160000 127.360000 ;
      RECT 547.100000 126.280000 548.960000 127.030000 ;
      RECT 506.620000 126.280000 545.300000 127.360000 ;
      RECT 461.620000 126.280000 504.820000 127.360000 ;
      RECT 416.620000 126.280000 459.820000 127.360000 ;
      RECT 371.620000 126.280000 414.820000 127.360000 ;
      RECT 326.620000 126.280000 369.820000 127.360000 ;
      RECT 281.620000 126.280000 324.820000 127.360000 ;
      RECT 236.620000 126.280000 279.820000 127.360000 ;
      RECT 191.620000 126.280000 234.820000 127.360000 ;
      RECT 146.620000 126.280000 189.820000 127.360000 ;
      RECT 101.620000 126.280000 144.820000 127.360000 ;
      RECT 56.620000 126.280000 99.820000 127.360000 ;
      RECT 11.620000 126.280000 54.820000 127.360000 ;
      RECT 4.860000 126.280000 9.655000 127.360000 ;
      RECT 0.000000 126.280000 3.060000 127.360000 ;
      RECT 0.000000 126.050000 548.960000 126.280000 ;
      RECT 0.000000 124.640000 550.160000 126.050000 ;
      RECT 544.900000 123.560000 550.160000 124.640000 ;
      RECT 508.620000 123.560000 543.100000 124.640000 ;
      RECT 463.620000 123.560000 506.820000 124.640000 ;
      RECT 418.620000 123.560000 461.820000 124.640000 ;
      RECT 373.620000 123.560000 416.820000 124.640000 ;
      RECT 328.620000 123.560000 371.820000 124.640000 ;
      RECT 283.620000 123.560000 326.820000 124.640000 ;
      RECT 238.620000 123.560000 281.820000 124.640000 ;
      RECT 193.620000 123.560000 236.820000 124.640000 ;
      RECT 148.620000 123.560000 191.820000 124.640000 ;
      RECT 103.620000 123.560000 146.820000 124.640000 ;
      RECT 58.620000 123.560000 101.820000 124.640000 ;
      RECT 13.620000 123.560000 56.820000 124.640000 ;
      RECT 7.060000 123.560000 11.820000 124.640000 ;
      RECT 0.000000 123.560000 5.260000 124.640000 ;
      RECT 0.000000 123.370000 550.160000 123.560000 ;
      RECT 0.000000 122.390000 548.960000 123.370000 ;
      RECT 0.000000 121.920000 550.160000 122.390000 ;
      RECT 547.100000 120.840000 550.160000 121.920000 ;
      RECT 506.620000 120.840000 545.300000 121.920000 ;
      RECT 461.620000 120.840000 504.820000 121.920000 ;
      RECT 416.620000 120.840000 459.820000 121.920000 ;
      RECT 371.620000 120.840000 414.820000 121.920000 ;
      RECT 326.620000 120.840000 369.820000 121.920000 ;
      RECT 281.620000 120.840000 324.820000 121.920000 ;
      RECT 236.620000 120.840000 279.820000 121.920000 ;
      RECT 191.620000 120.840000 234.820000 121.920000 ;
      RECT 146.620000 120.840000 189.820000 121.920000 ;
      RECT 101.620000 120.840000 144.820000 121.920000 ;
      RECT 56.620000 120.840000 99.820000 121.920000 ;
      RECT 11.620000 120.840000 54.820000 121.920000 ;
      RECT 4.860000 120.840000 9.655000 121.920000 ;
      RECT 0.000000 120.840000 3.060000 121.920000 ;
      RECT 0.000000 120.320000 550.160000 120.840000 ;
      RECT 0.000000 119.340000 548.960000 120.320000 ;
      RECT 0.000000 119.200000 550.160000 119.340000 ;
      RECT 544.900000 118.120000 550.160000 119.200000 ;
      RECT 508.620000 118.120000 543.100000 119.200000 ;
      RECT 463.620000 118.120000 506.820000 119.200000 ;
      RECT 418.620000 118.120000 461.820000 119.200000 ;
      RECT 373.620000 118.120000 416.820000 119.200000 ;
      RECT 328.620000 118.120000 371.820000 119.200000 ;
      RECT 283.620000 118.120000 326.820000 119.200000 ;
      RECT 238.620000 118.120000 281.820000 119.200000 ;
      RECT 193.620000 118.120000 236.820000 119.200000 ;
      RECT 148.620000 118.120000 191.820000 119.200000 ;
      RECT 103.620000 118.120000 146.820000 119.200000 ;
      RECT 58.620000 118.120000 101.820000 119.200000 ;
      RECT 13.620000 118.120000 56.820000 119.200000 ;
      RECT 7.060000 118.120000 11.820000 119.200000 ;
      RECT 0.000000 118.120000 5.260000 119.200000 ;
      RECT 0.000000 117.270000 550.160000 118.120000 ;
      RECT 0.000000 116.480000 548.960000 117.270000 ;
      RECT 547.100000 116.290000 548.960000 116.480000 ;
      RECT 547.100000 115.400000 550.160000 116.290000 ;
      RECT 506.620000 115.400000 545.300000 116.480000 ;
      RECT 461.620000 115.400000 504.820000 116.480000 ;
      RECT 416.620000 115.400000 459.820000 116.480000 ;
      RECT 371.620000 115.400000 414.820000 116.480000 ;
      RECT 326.620000 115.400000 369.820000 116.480000 ;
      RECT 281.620000 115.400000 324.820000 116.480000 ;
      RECT 236.620000 115.400000 279.820000 116.480000 ;
      RECT 191.620000 115.400000 234.820000 116.480000 ;
      RECT 146.620000 115.400000 189.820000 116.480000 ;
      RECT 101.620000 115.400000 144.820000 116.480000 ;
      RECT 56.620000 115.400000 99.820000 116.480000 ;
      RECT 11.620000 115.400000 54.820000 116.480000 ;
      RECT 4.860000 115.400000 9.655000 116.480000 ;
      RECT 0.000000 115.400000 3.060000 116.480000 ;
      RECT 0.000000 114.220000 550.160000 115.400000 ;
      RECT 0.000000 113.760000 548.960000 114.220000 ;
      RECT 544.900000 113.240000 548.960000 113.760000 ;
      RECT 544.900000 112.680000 550.160000 113.240000 ;
      RECT 508.620000 112.680000 543.100000 113.760000 ;
      RECT 463.620000 112.680000 506.820000 113.760000 ;
      RECT 418.620000 112.680000 461.820000 113.760000 ;
      RECT 373.620000 112.680000 416.820000 113.760000 ;
      RECT 328.620000 112.680000 371.820000 113.760000 ;
      RECT 283.620000 112.680000 326.820000 113.760000 ;
      RECT 238.620000 112.680000 281.820000 113.760000 ;
      RECT 193.620000 112.680000 236.820000 113.760000 ;
      RECT 148.620000 112.680000 191.820000 113.760000 ;
      RECT 103.620000 112.680000 146.820000 113.760000 ;
      RECT 58.620000 112.680000 101.820000 113.760000 ;
      RECT 13.620000 112.680000 56.820000 113.760000 ;
      RECT 7.060000 112.680000 11.820000 113.760000 ;
      RECT 0.000000 112.680000 5.260000 113.760000 ;
      RECT 0.000000 111.170000 550.160000 112.680000 ;
      RECT 0.000000 111.040000 548.960000 111.170000 ;
      RECT 547.100000 110.190000 548.960000 111.040000 ;
      RECT 547.100000 109.960000 550.160000 110.190000 ;
      RECT 506.620000 109.960000 545.300000 111.040000 ;
      RECT 461.620000 109.960000 504.820000 111.040000 ;
      RECT 416.620000 109.960000 459.820000 111.040000 ;
      RECT 371.620000 109.960000 414.820000 111.040000 ;
      RECT 326.620000 109.960000 369.820000 111.040000 ;
      RECT 281.620000 109.960000 324.820000 111.040000 ;
      RECT 236.620000 109.960000 279.820000 111.040000 ;
      RECT 191.620000 109.960000 234.820000 111.040000 ;
      RECT 146.620000 109.960000 189.820000 111.040000 ;
      RECT 101.620000 109.960000 144.820000 111.040000 ;
      RECT 56.620000 109.960000 99.820000 111.040000 ;
      RECT 11.620000 109.960000 54.820000 111.040000 ;
      RECT 4.860000 109.960000 9.655000 111.040000 ;
      RECT 0.000000 109.960000 3.060000 111.040000 ;
      RECT 0.000000 108.320000 550.160000 109.960000 ;
      RECT 544.900000 108.120000 550.160000 108.320000 ;
      RECT 544.900000 107.240000 548.960000 108.120000 ;
      RECT 508.620000 107.240000 543.100000 108.320000 ;
      RECT 463.620000 107.240000 506.820000 108.320000 ;
      RECT 418.620000 107.240000 461.820000 108.320000 ;
      RECT 373.620000 107.240000 416.820000 108.320000 ;
      RECT 328.620000 107.240000 371.820000 108.320000 ;
      RECT 283.620000 107.240000 326.820000 108.320000 ;
      RECT 238.620000 107.240000 281.820000 108.320000 ;
      RECT 193.620000 107.240000 236.820000 108.320000 ;
      RECT 148.620000 107.240000 191.820000 108.320000 ;
      RECT 103.620000 107.240000 146.820000 108.320000 ;
      RECT 58.620000 107.240000 101.820000 108.320000 ;
      RECT 13.620000 107.240000 56.820000 108.320000 ;
      RECT 7.060000 107.240000 11.820000 108.320000 ;
      RECT 0.000000 107.240000 5.260000 108.320000 ;
      RECT 0.000000 107.140000 548.960000 107.240000 ;
      RECT 0.000000 105.600000 550.160000 107.140000 ;
      RECT 547.100000 105.070000 550.160000 105.600000 ;
      RECT 547.100000 104.520000 548.960000 105.070000 ;
      RECT 506.620000 104.520000 545.300000 105.600000 ;
      RECT 461.620000 104.520000 504.820000 105.600000 ;
      RECT 416.620000 104.520000 459.820000 105.600000 ;
      RECT 371.620000 104.520000 414.820000 105.600000 ;
      RECT 326.620000 104.520000 369.820000 105.600000 ;
      RECT 281.620000 104.520000 324.820000 105.600000 ;
      RECT 236.620000 104.520000 279.820000 105.600000 ;
      RECT 191.620000 104.520000 234.820000 105.600000 ;
      RECT 146.620000 104.520000 189.820000 105.600000 ;
      RECT 101.620000 104.520000 144.820000 105.600000 ;
      RECT 56.620000 104.520000 99.820000 105.600000 ;
      RECT 11.620000 104.520000 54.820000 105.600000 ;
      RECT 4.860000 104.520000 9.655000 105.600000 ;
      RECT 0.000000 104.520000 3.060000 105.600000 ;
      RECT 0.000000 104.090000 548.960000 104.520000 ;
      RECT 0.000000 102.880000 550.160000 104.090000 ;
      RECT 544.900000 101.800000 550.160000 102.880000 ;
      RECT 508.620000 101.800000 543.100000 102.880000 ;
      RECT 463.620000 101.800000 506.820000 102.880000 ;
      RECT 418.620000 101.800000 461.820000 102.880000 ;
      RECT 373.620000 101.800000 416.820000 102.880000 ;
      RECT 328.620000 101.800000 371.820000 102.880000 ;
      RECT 283.620000 101.800000 326.820000 102.880000 ;
      RECT 238.620000 101.800000 281.820000 102.880000 ;
      RECT 193.620000 101.800000 236.820000 102.880000 ;
      RECT 148.620000 101.800000 191.820000 102.880000 ;
      RECT 103.620000 101.800000 146.820000 102.880000 ;
      RECT 58.620000 101.800000 101.820000 102.880000 ;
      RECT 13.620000 101.800000 56.820000 102.880000 ;
      RECT 7.060000 101.800000 11.820000 102.880000 ;
      RECT 0.000000 101.800000 5.260000 102.880000 ;
      RECT 0.000000 101.410000 550.160000 101.800000 ;
      RECT 0.000000 100.430000 548.960000 101.410000 ;
      RECT 0.000000 100.160000 550.160000 100.430000 ;
      RECT 547.100000 99.080000 550.160000 100.160000 ;
      RECT 506.620000 99.080000 545.300000 100.160000 ;
      RECT 461.620000 99.080000 504.820000 100.160000 ;
      RECT 416.620000 99.080000 459.820000 100.160000 ;
      RECT 371.620000 99.080000 414.820000 100.160000 ;
      RECT 326.620000 99.080000 369.820000 100.160000 ;
      RECT 281.620000 99.080000 324.820000 100.160000 ;
      RECT 236.620000 99.080000 279.820000 100.160000 ;
      RECT 191.620000 99.080000 234.820000 100.160000 ;
      RECT 146.620000 99.080000 189.820000 100.160000 ;
      RECT 101.620000 99.080000 144.820000 100.160000 ;
      RECT 56.620000 99.080000 99.820000 100.160000 ;
      RECT 11.620000 99.080000 54.820000 100.160000 ;
      RECT 4.860000 99.080000 9.655000 100.160000 ;
      RECT 0.000000 99.080000 3.060000 100.160000 ;
      RECT 0.000000 98.360000 550.160000 99.080000 ;
      RECT 0.000000 97.440000 548.960000 98.360000 ;
      RECT 544.900000 97.380000 548.960000 97.440000 ;
      RECT 544.900000 96.360000 550.160000 97.380000 ;
      RECT 508.620000 96.360000 543.100000 97.440000 ;
      RECT 463.620000 96.360000 506.820000 97.440000 ;
      RECT 418.620000 96.360000 461.820000 97.440000 ;
      RECT 373.620000 96.360000 416.820000 97.440000 ;
      RECT 328.620000 96.360000 371.820000 97.440000 ;
      RECT 283.620000 96.360000 326.820000 97.440000 ;
      RECT 238.620000 96.360000 281.820000 97.440000 ;
      RECT 193.620000 96.360000 236.820000 97.440000 ;
      RECT 148.620000 96.360000 191.820000 97.440000 ;
      RECT 103.620000 96.360000 146.820000 97.440000 ;
      RECT 58.620000 96.360000 101.820000 97.440000 ;
      RECT 13.620000 96.360000 56.820000 97.440000 ;
      RECT 7.060000 96.360000 11.820000 97.440000 ;
      RECT 0.000000 96.360000 5.260000 97.440000 ;
      RECT 0.000000 95.310000 550.160000 96.360000 ;
      RECT 0.000000 94.720000 548.960000 95.310000 ;
      RECT 547.100000 94.330000 548.960000 94.720000 ;
      RECT 547.100000 93.640000 550.160000 94.330000 ;
      RECT 506.620000 93.640000 545.300000 94.720000 ;
      RECT 461.620000 93.640000 504.820000 94.720000 ;
      RECT 416.620000 93.640000 459.820000 94.720000 ;
      RECT 371.620000 93.640000 414.820000 94.720000 ;
      RECT 326.620000 93.640000 369.820000 94.720000 ;
      RECT 281.620000 93.640000 324.820000 94.720000 ;
      RECT 236.620000 93.640000 279.820000 94.720000 ;
      RECT 191.620000 93.640000 234.820000 94.720000 ;
      RECT 146.620000 93.640000 189.820000 94.720000 ;
      RECT 101.620000 93.640000 144.820000 94.720000 ;
      RECT 56.620000 93.640000 99.820000 94.720000 ;
      RECT 11.620000 93.640000 54.820000 94.720000 ;
      RECT 4.860000 93.640000 9.655000 94.720000 ;
      RECT 0.000000 93.640000 3.060000 94.720000 ;
      RECT 0.000000 92.260000 550.160000 93.640000 ;
      RECT 0.000000 92.000000 548.960000 92.260000 ;
      RECT 544.900000 91.280000 548.960000 92.000000 ;
      RECT 544.900000 90.920000 550.160000 91.280000 ;
      RECT 508.620000 90.920000 543.100000 92.000000 ;
      RECT 463.620000 90.920000 506.820000 92.000000 ;
      RECT 418.620000 90.920000 461.820000 92.000000 ;
      RECT 373.620000 90.920000 416.820000 92.000000 ;
      RECT 328.620000 90.920000 371.820000 92.000000 ;
      RECT 283.620000 90.920000 326.820000 92.000000 ;
      RECT 238.620000 90.920000 281.820000 92.000000 ;
      RECT 193.620000 90.920000 236.820000 92.000000 ;
      RECT 148.620000 90.920000 191.820000 92.000000 ;
      RECT 103.620000 90.920000 146.820000 92.000000 ;
      RECT 58.620000 90.920000 101.820000 92.000000 ;
      RECT 13.620000 90.920000 56.820000 92.000000 ;
      RECT 7.060000 90.920000 11.820000 92.000000 ;
      RECT 0.000000 90.920000 5.260000 92.000000 ;
      RECT 0.000000 89.280000 550.160000 90.920000 ;
      RECT 547.100000 89.210000 550.160000 89.280000 ;
      RECT 547.100000 88.230000 548.960000 89.210000 ;
      RECT 547.100000 88.200000 550.160000 88.230000 ;
      RECT 506.620000 88.200000 545.300000 89.280000 ;
      RECT 461.620000 88.200000 504.820000 89.280000 ;
      RECT 416.620000 88.200000 459.820000 89.280000 ;
      RECT 371.620000 88.200000 414.820000 89.280000 ;
      RECT 326.620000 88.200000 369.820000 89.280000 ;
      RECT 281.620000 88.200000 324.820000 89.280000 ;
      RECT 236.620000 88.200000 279.820000 89.280000 ;
      RECT 191.620000 88.200000 234.820000 89.280000 ;
      RECT 146.620000 88.200000 189.820000 89.280000 ;
      RECT 101.620000 88.200000 144.820000 89.280000 ;
      RECT 56.620000 88.200000 99.820000 89.280000 ;
      RECT 11.620000 88.200000 54.820000 89.280000 ;
      RECT 4.860000 88.200000 9.655000 89.280000 ;
      RECT 0.000000 88.200000 3.060000 89.280000 ;
      RECT 0.000000 86.560000 550.160000 88.200000 ;
      RECT 544.900000 86.160000 550.160000 86.560000 ;
      RECT 544.900000 85.480000 548.960000 86.160000 ;
      RECT 508.620000 85.480000 543.100000 86.560000 ;
      RECT 463.620000 85.480000 506.820000 86.560000 ;
      RECT 418.620000 85.480000 461.820000 86.560000 ;
      RECT 373.620000 85.480000 416.820000 86.560000 ;
      RECT 328.620000 85.480000 371.820000 86.560000 ;
      RECT 283.620000 85.480000 326.820000 86.560000 ;
      RECT 238.620000 85.480000 281.820000 86.560000 ;
      RECT 193.620000 85.480000 236.820000 86.560000 ;
      RECT 148.620000 85.480000 191.820000 86.560000 ;
      RECT 103.620000 85.480000 146.820000 86.560000 ;
      RECT 58.620000 85.480000 101.820000 86.560000 ;
      RECT 13.620000 85.480000 56.820000 86.560000 ;
      RECT 7.060000 85.480000 11.820000 86.560000 ;
      RECT 0.000000 85.480000 5.260000 86.560000 ;
      RECT 0.000000 85.180000 548.960000 85.480000 ;
      RECT 0.000000 83.840000 550.160000 85.180000 ;
      RECT 547.100000 82.760000 550.160000 83.840000 ;
      RECT 506.620000 82.760000 545.300000 83.840000 ;
      RECT 461.620000 82.760000 504.820000 83.840000 ;
      RECT 416.620000 82.760000 459.820000 83.840000 ;
      RECT 371.620000 82.760000 414.820000 83.840000 ;
      RECT 326.620000 82.760000 369.820000 83.840000 ;
      RECT 281.620000 82.760000 324.820000 83.840000 ;
      RECT 236.620000 82.760000 279.820000 83.840000 ;
      RECT 191.620000 82.760000 234.820000 83.840000 ;
      RECT 146.620000 82.760000 189.820000 83.840000 ;
      RECT 101.620000 82.760000 144.820000 83.840000 ;
      RECT 56.620000 82.760000 99.820000 83.840000 ;
      RECT 11.620000 82.760000 54.820000 83.840000 ;
      RECT 4.860000 82.760000 9.655000 83.840000 ;
      RECT 0.000000 82.760000 3.060000 83.840000 ;
      RECT 0.000000 82.500000 550.160000 82.760000 ;
      RECT 0.000000 81.520000 548.960000 82.500000 ;
      RECT 0.000000 81.120000 550.160000 81.520000 ;
      RECT 544.900000 80.040000 550.160000 81.120000 ;
      RECT 508.620000 80.040000 543.100000 81.120000 ;
      RECT 463.620000 80.040000 506.820000 81.120000 ;
      RECT 418.620000 80.040000 461.820000 81.120000 ;
      RECT 373.620000 80.040000 416.820000 81.120000 ;
      RECT 328.620000 80.040000 371.820000 81.120000 ;
      RECT 283.620000 80.040000 326.820000 81.120000 ;
      RECT 238.620000 80.040000 281.820000 81.120000 ;
      RECT 193.620000 80.040000 236.820000 81.120000 ;
      RECT 148.620000 80.040000 191.820000 81.120000 ;
      RECT 103.620000 80.040000 146.820000 81.120000 ;
      RECT 58.620000 80.040000 101.820000 81.120000 ;
      RECT 13.620000 80.040000 56.820000 81.120000 ;
      RECT 7.060000 80.040000 11.820000 81.120000 ;
      RECT 0.000000 80.040000 5.260000 81.120000 ;
      RECT 0.000000 79.450000 550.160000 80.040000 ;
      RECT 0.000000 78.470000 548.960000 79.450000 ;
      RECT 0.000000 78.400000 550.160000 78.470000 ;
      RECT 547.100000 77.320000 550.160000 78.400000 ;
      RECT 506.620000 77.320000 545.300000 78.400000 ;
      RECT 461.620000 77.320000 504.820000 78.400000 ;
      RECT 416.620000 77.320000 459.820000 78.400000 ;
      RECT 371.620000 77.320000 414.820000 78.400000 ;
      RECT 326.620000 77.320000 369.820000 78.400000 ;
      RECT 281.620000 77.320000 324.820000 78.400000 ;
      RECT 236.620000 77.320000 279.820000 78.400000 ;
      RECT 191.620000 77.320000 234.820000 78.400000 ;
      RECT 146.620000 77.320000 189.820000 78.400000 ;
      RECT 101.620000 77.320000 144.820000 78.400000 ;
      RECT 56.620000 77.320000 99.820000 78.400000 ;
      RECT 11.620000 77.320000 54.820000 78.400000 ;
      RECT 4.860000 77.320000 9.655000 78.400000 ;
      RECT 0.000000 77.320000 3.060000 78.400000 ;
      RECT 0.000000 76.400000 550.160000 77.320000 ;
      RECT 0.000000 75.680000 548.960000 76.400000 ;
      RECT 544.900000 75.420000 548.960000 75.680000 ;
      RECT 544.900000 74.600000 550.160000 75.420000 ;
      RECT 508.620000 74.600000 543.100000 75.680000 ;
      RECT 463.620000 74.600000 506.820000 75.680000 ;
      RECT 418.620000 74.600000 461.820000 75.680000 ;
      RECT 373.620000 74.600000 416.820000 75.680000 ;
      RECT 328.620000 74.600000 371.820000 75.680000 ;
      RECT 283.620000 74.600000 326.820000 75.680000 ;
      RECT 238.620000 74.600000 281.820000 75.680000 ;
      RECT 193.620000 74.600000 236.820000 75.680000 ;
      RECT 148.620000 74.600000 191.820000 75.680000 ;
      RECT 103.620000 74.600000 146.820000 75.680000 ;
      RECT 58.620000 74.600000 101.820000 75.680000 ;
      RECT 13.620000 74.600000 56.820000 75.680000 ;
      RECT 7.060000 74.600000 11.820000 75.680000 ;
      RECT 0.000000 74.600000 5.260000 75.680000 ;
      RECT 0.000000 73.350000 550.160000 74.600000 ;
      RECT 0.000000 72.960000 548.960000 73.350000 ;
      RECT 547.100000 72.370000 548.960000 72.960000 ;
      RECT 547.100000 71.880000 550.160000 72.370000 ;
      RECT 506.620000 71.880000 545.300000 72.960000 ;
      RECT 461.620000 71.880000 504.820000 72.960000 ;
      RECT 416.620000 71.880000 459.820000 72.960000 ;
      RECT 371.620000 71.880000 414.820000 72.960000 ;
      RECT 326.620000 71.880000 369.820000 72.960000 ;
      RECT 281.620000 71.880000 324.820000 72.960000 ;
      RECT 236.620000 71.880000 279.820000 72.960000 ;
      RECT 191.620000 71.880000 234.820000 72.960000 ;
      RECT 146.620000 71.880000 189.820000 72.960000 ;
      RECT 101.620000 71.880000 144.820000 72.960000 ;
      RECT 56.620000 71.880000 99.820000 72.960000 ;
      RECT 11.620000 71.880000 54.820000 72.960000 ;
      RECT 4.860000 71.880000 9.655000 72.960000 ;
      RECT 0.000000 71.880000 3.060000 72.960000 ;
      RECT 0.000000 70.300000 550.160000 71.880000 ;
      RECT 0.000000 70.240000 548.960000 70.300000 ;
      RECT 544.900000 69.320000 548.960000 70.240000 ;
      RECT 544.900000 69.160000 550.160000 69.320000 ;
      RECT 508.620000 69.160000 543.100000 70.240000 ;
      RECT 463.620000 69.160000 506.820000 70.240000 ;
      RECT 418.620000 69.160000 461.820000 70.240000 ;
      RECT 373.620000 69.160000 416.820000 70.240000 ;
      RECT 328.620000 69.160000 371.820000 70.240000 ;
      RECT 283.620000 69.160000 326.820000 70.240000 ;
      RECT 238.620000 69.160000 281.820000 70.240000 ;
      RECT 193.620000 69.160000 236.820000 70.240000 ;
      RECT 148.620000 69.160000 191.820000 70.240000 ;
      RECT 103.620000 69.160000 146.820000 70.240000 ;
      RECT 58.620000 69.160000 101.820000 70.240000 ;
      RECT 13.620000 69.160000 56.820000 70.240000 ;
      RECT 7.060000 69.160000 11.820000 70.240000 ;
      RECT 0.000000 69.160000 5.260000 70.240000 ;
      RECT 0.000000 67.520000 550.160000 69.160000 ;
      RECT 547.100000 67.250000 550.160000 67.520000 ;
      RECT 547.100000 66.440000 548.960000 67.250000 ;
      RECT 506.620000 66.440000 545.300000 67.520000 ;
      RECT 461.620000 66.440000 504.820000 67.520000 ;
      RECT 416.620000 66.440000 459.820000 67.520000 ;
      RECT 371.620000 66.440000 414.820000 67.520000 ;
      RECT 326.620000 66.440000 369.820000 67.520000 ;
      RECT 281.620000 66.440000 324.820000 67.520000 ;
      RECT 236.620000 66.440000 279.820000 67.520000 ;
      RECT 191.620000 66.440000 234.820000 67.520000 ;
      RECT 146.620000 66.440000 189.820000 67.520000 ;
      RECT 101.620000 66.440000 144.820000 67.520000 ;
      RECT 56.620000 66.440000 99.820000 67.520000 ;
      RECT 11.620000 66.440000 54.820000 67.520000 ;
      RECT 4.860000 66.440000 9.655000 67.520000 ;
      RECT 0.000000 66.440000 3.060000 67.520000 ;
      RECT 0.000000 66.270000 548.960000 66.440000 ;
      RECT 0.000000 64.800000 550.160000 66.270000 ;
      RECT 544.900000 63.720000 550.160000 64.800000 ;
      RECT 508.620000 63.720000 543.100000 64.800000 ;
      RECT 463.620000 63.720000 506.820000 64.800000 ;
      RECT 418.620000 63.720000 461.820000 64.800000 ;
      RECT 373.620000 63.720000 416.820000 64.800000 ;
      RECT 328.620000 63.720000 371.820000 64.800000 ;
      RECT 283.620000 63.720000 326.820000 64.800000 ;
      RECT 238.620000 63.720000 281.820000 64.800000 ;
      RECT 193.620000 63.720000 236.820000 64.800000 ;
      RECT 148.620000 63.720000 191.820000 64.800000 ;
      RECT 103.620000 63.720000 146.820000 64.800000 ;
      RECT 58.620000 63.720000 101.820000 64.800000 ;
      RECT 13.620000 63.720000 56.820000 64.800000 ;
      RECT 7.060000 63.720000 11.820000 64.800000 ;
      RECT 0.000000 63.720000 5.260000 64.800000 ;
      RECT 0.000000 63.590000 550.160000 63.720000 ;
      RECT 0.000000 62.610000 548.960000 63.590000 ;
      RECT 0.000000 62.080000 550.160000 62.610000 ;
      RECT 547.100000 61.000000 550.160000 62.080000 ;
      RECT 506.620000 61.000000 545.300000 62.080000 ;
      RECT 461.620000 61.000000 504.820000 62.080000 ;
      RECT 416.620000 61.000000 459.820000 62.080000 ;
      RECT 371.620000 61.000000 414.820000 62.080000 ;
      RECT 326.620000 61.000000 369.820000 62.080000 ;
      RECT 281.620000 61.000000 324.820000 62.080000 ;
      RECT 236.620000 61.000000 279.820000 62.080000 ;
      RECT 191.620000 61.000000 234.820000 62.080000 ;
      RECT 146.620000 61.000000 189.820000 62.080000 ;
      RECT 101.620000 61.000000 144.820000 62.080000 ;
      RECT 56.620000 61.000000 99.820000 62.080000 ;
      RECT 11.620000 61.000000 54.820000 62.080000 ;
      RECT 4.860000 61.000000 9.655000 62.080000 ;
      RECT 0.000000 61.000000 3.060000 62.080000 ;
      RECT 0.000000 60.540000 550.160000 61.000000 ;
      RECT 0.000000 59.560000 548.960000 60.540000 ;
      RECT 0.000000 59.360000 550.160000 59.560000 ;
      RECT 544.900000 58.280000 550.160000 59.360000 ;
      RECT 508.620000 58.280000 543.100000 59.360000 ;
      RECT 463.620000 58.280000 506.820000 59.360000 ;
      RECT 418.620000 58.280000 461.820000 59.360000 ;
      RECT 373.620000 58.280000 416.820000 59.360000 ;
      RECT 328.620000 58.280000 371.820000 59.360000 ;
      RECT 283.620000 58.280000 326.820000 59.360000 ;
      RECT 238.620000 58.280000 281.820000 59.360000 ;
      RECT 193.620000 58.280000 236.820000 59.360000 ;
      RECT 148.620000 58.280000 191.820000 59.360000 ;
      RECT 103.620000 58.280000 146.820000 59.360000 ;
      RECT 58.620000 58.280000 101.820000 59.360000 ;
      RECT 13.620000 58.280000 56.820000 59.360000 ;
      RECT 7.060000 58.280000 11.820000 59.360000 ;
      RECT 0.000000 58.280000 5.260000 59.360000 ;
      RECT 0.000000 57.490000 550.160000 58.280000 ;
      RECT 0.000000 56.640000 548.960000 57.490000 ;
      RECT 547.100000 56.510000 548.960000 56.640000 ;
      RECT 547.100000 55.560000 550.160000 56.510000 ;
      RECT 506.620000 55.560000 545.300000 56.640000 ;
      RECT 461.620000 55.560000 504.820000 56.640000 ;
      RECT 416.620000 55.560000 459.820000 56.640000 ;
      RECT 371.620000 55.560000 414.820000 56.640000 ;
      RECT 326.620000 55.560000 369.820000 56.640000 ;
      RECT 281.620000 55.560000 324.820000 56.640000 ;
      RECT 236.620000 55.560000 279.820000 56.640000 ;
      RECT 191.620000 55.560000 234.820000 56.640000 ;
      RECT 146.620000 55.560000 189.820000 56.640000 ;
      RECT 101.620000 55.560000 144.820000 56.640000 ;
      RECT 56.620000 55.560000 99.820000 56.640000 ;
      RECT 11.620000 55.560000 54.820000 56.640000 ;
      RECT 4.860000 55.560000 9.655000 56.640000 ;
      RECT 0.000000 55.560000 3.060000 56.640000 ;
      RECT 0.000000 54.440000 550.160000 55.560000 ;
      RECT 0.000000 53.920000 548.960000 54.440000 ;
      RECT 544.900000 53.460000 548.960000 53.920000 ;
      RECT 544.900000 52.840000 550.160000 53.460000 ;
      RECT 508.620000 52.840000 543.100000 53.920000 ;
      RECT 463.620000 52.840000 506.820000 53.920000 ;
      RECT 418.620000 52.840000 461.820000 53.920000 ;
      RECT 373.620000 52.840000 416.820000 53.920000 ;
      RECT 328.620000 52.840000 371.820000 53.920000 ;
      RECT 283.620000 52.840000 326.820000 53.920000 ;
      RECT 238.620000 52.840000 281.820000 53.920000 ;
      RECT 193.620000 52.840000 236.820000 53.920000 ;
      RECT 148.620000 52.840000 191.820000 53.920000 ;
      RECT 103.620000 52.840000 146.820000 53.920000 ;
      RECT 58.620000 52.840000 101.820000 53.920000 ;
      RECT 13.620000 52.840000 56.820000 53.920000 ;
      RECT 7.060000 52.840000 11.820000 53.920000 ;
      RECT 0.000000 52.840000 5.260000 53.920000 ;
      RECT 0.000000 51.390000 550.160000 52.840000 ;
      RECT 0.000000 51.200000 548.960000 51.390000 ;
      RECT 547.100000 50.410000 548.960000 51.200000 ;
      RECT 547.100000 50.120000 550.160000 50.410000 ;
      RECT 506.620000 50.120000 545.300000 51.200000 ;
      RECT 461.620000 50.120000 504.820000 51.200000 ;
      RECT 416.620000 50.120000 459.820000 51.200000 ;
      RECT 371.620000 50.120000 414.820000 51.200000 ;
      RECT 326.620000 50.120000 369.820000 51.200000 ;
      RECT 281.620000 50.120000 324.820000 51.200000 ;
      RECT 236.620000 50.120000 279.820000 51.200000 ;
      RECT 191.620000 50.120000 234.820000 51.200000 ;
      RECT 146.620000 50.120000 189.820000 51.200000 ;
      RECT 101.620000 50.120000 144.820000 51.200000 ;
      RECT 56.620000 50.120000 99.820000 51.200000 ;
      RECT 11.620000 50.120000 54.820000 51.200000 ;
      RECT 4.860000 50.120000 9.655000 51.200000 ;
      RECT 0.000000 50.120000 3.060000 51.200000 ;
      RECT 0.000000 48.480000 550.160000 50.120000 ;
      RECT 544.900000 47.730000 550.160000 48.480000 ;
      RECT 544.900000 47.400000 548.960000 47.730000 ;
      RECT 508.620000 47.400000 543.100000 48.480000 ;
      RECT 463.620000 47.400000 506.820000 48.480000 ;
      RECT 418.620000 47.400000 461.820000 48.480000 ;
      RECT 373.620000 47.400000 416.820000 48.480000 ;
      RECT 328.620000 47.400000 371.820000 48.480000 ;
      RECT 283.620000 47.400000 326.820000 48.480000 ;
      RECT 238.620000 47.400000 281.820000 48.480000 ;
      RECT 193.620000 47.400000 236.820000 48.480000 ;
      RECT 148.620000 47.400000 191.820000 48.480000 ;
      RECT 103.620000 47.400000 146.820000 48.480000 ;
      RECT 58.620000 47.400000 101.820000 48.480000 ;
      RECT 13.620000 47.400000 56.820000 48.480000 ;
      RECT 7.060000 47.400000 11.820000 48.480000 ;
      RECT 0.000000 47.400000 5.260000 48.480000 ;
      RECT 0.000000 46.750000 548.960000 47.400000 ;
      RECT 0.000000 45.760000 550.160000 46.750000 ;
      RECT 547.100000 44.680000 550.160000 45.760000 ;
      RECT 506.620000 44.680000 545.300000 45.760000 ;
      RECT 461.620000 44.680000 504.820000 45.760000 ;
      RECT 416.620000 44.680000 459.820000 45.760000 ;
      RECT 371.620000 44.680000 414.820000 45.760000 ;
      RECT 326.620000 44.680000 369.820000 45.760000 ;
      RECT 281.620000 44.680000 324.820000 45.760000 ;
      RECT 236.620000 44.680000 279.820000 45.760000 ;
      RECT 191.620000 44.680000 234.820000 45.760000 ;
      RECT 146.620000 44.680000 189.820000 45.760000 ;
      RECT 101.620000 44.680000 144.820000 45.760000 ;
      RECT 56.620000 44.680000 99.820000 45.760000 ;
      RECT 11.620000 44.680000 54.820000 45.760000 ;
      RECT 4.860000 44.680000 9.655000 45.760000 ;
      RECT 0.000000 44.680000 3.060000 45.760000 ;
      RECT 0.000000 43.700000 548.960000 44.680000 ;
      RECT 0.000000 43.040000 550.160000 43.700000 ;
      RECT 544.900000 41.960000 550.160000 43.040000 ;
      RECT 508.620000 41.960000 543.100000 43.040000 ;
      RECT 463.620000 41.960000 506.820000 43.040000 ;
      RECT 418.620000 41.960000 461.820000 43.040000 ;
      RECT 373.620000 41.960000 416.820000 43.040000 ;
      RECT 328.620000 41.960000 371.820000 43.040000 ;
      RECT 283.620000 41.960000 326.820000 43.040000 ;
      RECT 238.620000 41.960000 281.820000 43.040000 ;
      RECT 193.620000 41.960000 236.820000 43.040000 ;
      RECT 148.620000 41.960000 191.820000 43.040000 ;
      RECT 103.620000 41.960000 146.820000 43.040000 ;
      RECT 58.620000 41.960000 101.820000 43.040000 ;
      RECT 13.620000 41.960000 56.820000 43.040000 ;
      RECT 7.060000 41.960000 11.820000 43.040000 ;
      RECT 0.000000 41.960000 5.260000 43.040000 ;
      RECT 0.000000 41.630000 550.160000 41.960000 ;
      RECT 0.000000 40.650000 548.960000 41.630000 ;
      RECT 0.000000 40.320000 550.160000 40.650000 ;
      RECT 547.100000 39.240000 550.160000 40.320000 ;
      RECT 506.620000 39.240000 545.300000 40.320000 ;
      RECT 461.620000 39.240000 504.820000 40.320000 ;
      RECT 416.620000 39.240000 459.820000 40.320000 ;
      RECT 371.620000 39.240000 414.820000 40.320000 ;
      RECT 326.620000 39.240000 369.820000 40.320000 ;
      RECT 281.620000 39.240000 324.820000 40.320000 ;
      RECT 236.620000 39.240000 279.820000 40.320000 ;
      RECT 191.620000 39.240000 234.820000 40.320000 ;
      RECT 146.620000 39.240000 189.820000 40.320000 ;
      RECT 101.620000 39.240000 144.820000 40.320000 ;
      RECT 56.620000 39.240000 99.820000 40.320000 ;
      RECT 11.620000 39.240000 54.820000 40.320000 ;
      RECT 4.860000 39.240000 9.655000 40.320000 ;
      RECT 0.000000 39.240000 3.060000 40.320000 ;
      RECT 0.000000 38.580000 550.160000 39.240000 ;
      RECT 0.000000 37.600000 548.960000 38.580000 ;
      RECT 544.900000 36.520000 550.160000 37.600000 ;
      RECT 508.620000 36.520000 543.100000 37.600000 ;
      RECT 463.620000 36.520000 506.820000 37.600000 ;
      RECT 418.620000 36.520000 461.820000 37.600000 ;
      RECT 373.620000 36.520000 416.820000 37.600000 ;
      RECT 328.620000 36.520000 371.820000 37.600000 ;
      RECT 283.620000 36.520000 326.820000 37.600000 ;
      RECT 238.620000 36.520000 281.820000 37.600000 ;
      RECT 193.620000 36.520000 236.820000 37.600000 ;
      RECT 148.620000 36.520000 191.820000 37.600000 ;
      RECT 103.620000 36.520000 146.820000 37.600000 ;
      RECT 58.620000 36.520000 101.820000 37.600000 ;
      RECT 13.620000 36.520000 56.820000 37.600000 ;
      RECT 7.060000 36.520000 11.820000 37.600000 ;
      RECT 0.000000 36.520000 5.260000 37.600000 ;
      RECT 0.000000 35.530000 550.160000 36.520000 ;
      RECT 0.000000 34.880000 548.960000 35.530000 ;
      RECT 547.100000 34.550000 548.960000 34.880000 ;
      RECT 547.100000 33.800000 550.160000 34.550000 ;
      RECT 506.620000 33.800000 545.300000 34.880000 ;
      RECT 461.620000 33.800000 504.820000 34.880000 ;
      RECT 416.620000 33.800000 459.820000 34.880000 ;
      RECT 371.620000 33.800000 414.820000 34.880000 ;
      RECT 326.620000 33.800000 369.820000 34.880000 ;
      RECT 281.620000 33.800000 324.820000 34.880000 ;
      RECT 236.620000 33.800000 279.820000 34.880000 ;
      RECT 191.620000 33.800000 234.820000 34.880000 ;
      RECT 146.620000 33.800000 189.820000 34.880000 ;
      RECT 101.620000 33.800000 144.820000 34.880000 ;
      RECT 56.620000 33.800000 99.820000 34.880000 ;
      RECT 11.620000 33.800000 54.820000 34.880000 ;
      RECT 4.860000 33.800000 9.655000 34.880000 ;
      RECT 0.000000 33.800000 3.060000 34.880000 ;
      RECT 0.000000 32.480000 550.160000 33.800000 ;
      RECT 0.000000 32.160000 548.960000 32.480000 ;
      RECT 544.900000 31.500000 548.960000 32.160000 ;
      RECT 544.900000 31.080000 550.160000 31.500000 ;
      RECT 508.620000 31.080000 543.100000 32.160000 ;
      RECT 463.620000 31.080000 506.820000 32.160000 ;
      RECT 418.620000 31.080000 461.820000 32.160000 ;
      RECT 373.620000 31.080000 416.820000 32.160000 ;
      RECT 328.620000 31.080000 371.820000 32.160000 ;
      RECT 283.620000 31.080000 326.820000 32.160000 ;
      RECT 238.620000 31.080000 281.820000 32.160000 ;
      RECT 193.620000 31.080000 236.820000 32.160000 ;
      RECT 148.620000 31.080000 191.820000 32.160000 ;
      RECT 103.620000 31.080000 146.820000 32.160000 ;
      RECT 58.620000 31.080000 101.820000 32.160000 ;
      RECT 13.620000 31.080000 56.820000 32.160000 ;
      RECT 7.060000 31.080000 11.820000 32.160000 ;
      RECT 0.000000 31.080000 5.260000 32.160000 ;
      RECT 0.000000 29.440000 550.160000 31.080000 ;
      RECT 547.100000 29.430000 550.160000 29.440000 ;
      RECT 547.100000 28.450000 548.960000 29.430000 ;
      RECT 547.100000 28.360000 550.160000 28.450000 ;
      RECT 506.620000 28.360000 545.300000 29.440000 ;
      RECT 461.620000 28.360000 504.820000 29.440000 ;
      RECT 416.620000 28.360000 459.820000 29.440000 ;
      RECT 371.620000 28.360000 414.820000 29.440000 ;
      RECT 326.620000 28.360000 369.820000 29.440000 ;
      RECT 281.620000 28.360000 324.820000 29.440000 ;
      RECT 236.620000 28.360000 279.820000 29.440000 ;
      RECT 191.620000 28.360000 234.820000 29.440000 ;
      RECT 146.620000 28.360000 189.820000 29.440000 ;
      RECT 101.620000 28.360000 144.820000 29.440000 ;
      RECT 56.620000 28.360000 99.820000 29.440000 ;
      RECT 11.620000 28.360000 54.820000 29.440000 ;
      RECT 4.860000 28.360000 9.655000 29.440000 ;
      RECT 0.000000 28.360000 3.060000 29.440000 ;
      RECT 0.000000 26.720000 550.160000 28.360000 ;
      RECT 544.900000 25.770000 550.160000 26.720000 ;
      RECT 544.900000 25.640000 548.960000 25.770000 ;
      RECT 508.620000 25.640000 543.100000 26.720000 ;
      RECT 463.620000 25.640000 506.820000 26.720000 ;
      RECT 418.620000 25.640000 461.820000 26.720000 ;
      RECT 373.620000 25.640000 416.820000 26.720000 ;
      RECT 328.620000 25.640000 371.820000 26.720000 ;
      RECT 283.620000 25.640000 326.820000 26.720000 ;
      RECT 238.620000 25.640000 281.820000 26.720000 ;
      RECT 193.620000 25.640000 236.820000 26.720000 ;
      RECT 148.620000 25.640000 191.820000 26.720000 ;
      RECT 103.620000 25.640000 146.820000 26.720000 ;
      RECT 58.620000 25.640000 101.820000 26.720000 ;
      RECT 13.620000 25.640000 56.820000 26.720000 ;
      RECT 7.060000 25.640000 11.820000 26.720000 ;
      RECT 0.000000 25.640000 5.260000 26.720000 ;
      RECT 0.000000 24.790000 548.960000 25.640000 ;
      RECT 0.000000 24.000000 550.160000 24.790000 ;
      RECT 547.100000 22.920000 550.160000 24.000000 ;
      RECT 506.620000 22.920000 545.300000 24.000000 ;
      RECT 461.620000 22.920000 504.820000 24.000000 ;
      RECT 416.620000 22.920000 459.820000 24.000000 ;
      RECT 371.620000 22.920000 414.820000 24.000000 ;
      RECT 326.620000 22.920000 369.820000 24.000000 ;
      RECT 281.620000 22.920000 324.820000 24.000000 ;
      RECT 236.620000 22.920000 279.820000 24.000000 ;
      RECT 191.620000 22.920000 234.820000 24.000000 ;
      RECT 146.620000 22.920000 189.820000 24.000000 ;
      RECT 101.620000 22.920000 144.820000 24.000000 ;
      RECT 56.620000 22.920000 99.820000 24.000000 ;
      RECT 11.620000 22.920000 54.820000 24.000000 ;
      RECT 4.860000 22.920000 9.655000 24.000000 ;
      RECT 0.000000 22.920000 3.060000 24.000000 ;
      RECT 0.000000 22.720000 550.160000 22.920000 ;
      RECT 0.000000 21.740000 548.960000 22.720000 ;
      RECT 0.000000 21.280000 550.160000 21.740000 ;
      RECT 544.900000 20.200000 550.160000 21.280000 ;
      RECT 508.620000 20.200000 543.100000 21.280000 ;
      RECT 463.620000 20.200000 506.820000 21.280000 ;
      RECT 418.620000 20.200000 461.820000 21.280000 ;
      RECT 373.620000 20.200000 416.820000 21.280000 ;
      RECT 328.620000 20.200000 371.820000 21.280000 ;
      RECT 283.620000 20.200000 326.820000 21.280000 ;
      RECT 238.620000 20.200000 281.820000 21.280000 ;
      RECT 193.620000 20.200000 236.820000 21.280000 ;
      RECT 148.620000 20.200000 191.820000 21.280000 ;
      RECT 103.620000 20.200000 146.820000 21.280000 ;
      RECT 58.620000 20.200000 101.820000 21.280000 ;
      RECT 13.620000 20.200000 56.820000 21.280000 ;
      RECT 7.060000 20.200000 11.820000 21.280000 ;
      RECT 0.000000 20.200000 5.260000 21.280000 ;
      RECT 0.000000 19.670000 550.160000 20.200000 ;
      RECT 0.000000 18.690000 548.960000 19.670000 ;
      RECT 0.000000 18.560000 550.160000 18.690000 ;
      RECT 547.100000 17.480000 550.160000 18.560000 ;
      RECT 506.620000 17.480000 545.300000 18.560000 ;
      RECT 461.620000 17.480000 504.820000 18.560000 ;
      RECT 416.620000 17.480000 459.820000 18.560000 ;
      RECT 371.620000 17.480000 414.820000 18.560000 ;
      RECT 326.620000 17.480000 369.820000 18.560000 ;
      RECT 281.620000 17.480000 324.820000 18.560000 ;
      RECT 236.620000 17.480000 279.820000 18.560000 ;
      RECT 191.620000 17.480000 234.820000 18.560000 ;
      RECT 146.620000 17.480000 189.820000 18.560000 ;
      RECT 101.620000 17.480000 144.820000 18.560000 ;
      RECT 56.620000 17.480000 99.820000 18.560000 ;
      RECT 11.620000 17.480000 54.820000 18.560000 ;
      RECT 4.860000 17.480000 9.655000 18.560000 ;
      RECT 0.000000 17.480000 3.060000 18.560000 ;
      RECT 0.000000 16.620000 550.160000 17.480000 ;
      RECT 0.000000 15.840000 548.960000 16.620000 ;
      RECT 544.900000 15.640000 548.960000 15.840000 ;
      RECT 544.900000 14.760000 550.160000 15.640000 ;
      RECT 508.620000 14.760000 543.100000 15.840000 ;
      RECT 463.620000 14.760000 506.820000 15.840000 ;
      RECT 418.620000 14.760000 461.820000 15.840000 ;
      RECT 373.620000 14.760000 416.820000 15.840000 ;
      RECT 328.620000 14.760000 371.820000 15.840000 ;
      RECT 283.620000 14.760000 326.820000 15.840000 ;
      RECT 238.620000 14.760000 281.820000 15.840000 ;
      RECT 193.620000 14.760000 236.820000 15.840000 ;
      RECT 148.620000 14.760000 191.820000 15.840000 ;
      RECT 103.620000 14.760000 146.820000 15.840000 ;
      RECT 58.620000 14.760000 101.820000 15.840000 ;
      RECT 13.620000 14.760000 56.820000 15.840000 ;
      RECT 7.060000 14.760000 11.820000 15.840000 ;
      RECT 0.000000 14.760000 5.260000 15.840000 ;
      RECT 0.000000 13.570000 550.160000 14.760000 ;
      RECT 0.000000 13.120000 548.960000 13.570000 ;
      RECT 547.100000 12.590000 548.960000 13.120000 ;
      RECT 547.100000 12.040000 550.160000 12.590000 ;
      RECT 506.620000 12.040000 545.300000 13.120000 ;
      RECT 461.620000 12.040000 504.820000 13.120000 ;
      RECT 416.620000 12.040000 459.820000 13.120000 ;
      RECT 371.620000 12.040000 414.820000 13.120000 ;
      RECT 326.620000 12.040000 369.820000 13.120000 ;
      RECT 281.620000 12.040000 324.820000 13.120000 ;
      RECT 236.620000 12.040000 279.820000 13.120000 ;
      RECT 191.620000 12.040000 234.820000 13.120000 ;
      RECT 146.620000 12.040000 189.820000 13.120000 ;
      RECT 101.620000 12.040000 144.820000 13.120000 ;
      RECT 56.620000 12.040000 99.820000 13.120000 ;
      RECT 11.620000 12.040000 54.820000 13.120000 ;
      RECT 4.860000 12.040000 9.655000 13.120000 ;
      RECT 0.000000 12.040000 3.060000 13.120000 ;
      RECT 0.000000 10.520000 550.160000 12.040000 ;
      RECT 0.000000 10.400000 548.960000 10.520000 ;
      RECT 544.900000 9.540000 548.960000 10.400000 ;
      RECT 544.900000 9.320000 550.160000 9.540000 ;
      RECT 508.620000 9.320000 543.100000 10.400000 ;
      RECT 463.620000 9.320000 506.820000 10.400000 ;
      RECT 418.620000 9.320000 461.820000 10.400000 ;
      RECT 373.620000 9.320000 416.820000 10.400000 ;
      RECT 328.620000 9.320000 371.820000 10.400000 ;
      RECT 283.620000 9.320000 326.820000 10.400000 ;
      RECT 238.620000 9.320000 281.820000 10.400000 ;
      RECT 193.620000 9.320000 236.820000 10.400000 ;
      RECT 148.620000 9.320000 191.820000 10.400000 ;
      RECT 103.620000 9.320000 146.820000 10.400000 ;
      RECT 58.620000 9.320000 101.820000 10.400000 ;
      RECT 13.620000 9.320000 56.820000 10.400000 ;
      RECT 7.060000 9.320000 11.820000 10.400000 ;
      RECT 0.000000 9.320000 5.260000 10.400000 ;
      RECT 0.000000 6.930000 550.160000 9.320000 ;
      RECT 0.000000 4.730000 550.160000 5.130000 ;
      RECT 0.000000 0.000000 550.160000 2.930000 ;
    LAYER met4 ;
      RECT 7.060000 545.660000 543.100000 549.780000 ;
      RECT 506.620000 543.460000 543.100000 545.660000 ;
      RECT 461.620000 543.460000 504.820000 545.660000 ;
      RECT 416.620000 543.460000 459.820000 545.660000 ;
      RECT 371.620000 543.460000 414.820000 545.660000 ;
      RECT 326.620000 543.460000 369.820000 545.660000 ;
      RECT 281.620000 543.460000 324.820000 545.660000 ;
      RECT 236.620000 543.460000 279.820000 545.660000 ;
      RECT 191.620000 543.460000 234.820000 545.660000 ;
      RECT 146.620000 543.460000 189.820000 545.660000 ;
      RECT 101.620000 543.460000 144.820000 545.660000 ;
      RECT 56.620000 543.460000 99.820000 545.660000 ;
      RECT 11.620000 543.460000 54.820000 545.660000 ;
      RECT 7.060000 535.360000 9.820000 545.660000 ;
      RECT 7.060000 534.280000 9.655000 535.360000 ;
      RECT 7.060000 529.920000 9.820000 534.280000 ;
      RECT 7.060000 528.840000 9.655000 529.920000 ;
      RECT 7.060000 524.480000 9.820000 528.840000 ;
      RECT 7.060000 523.400000 9.655000 524.480000 ;
      RECT 7.060000 519.040000 9.820000 523.400000 ;
      RECT 7.060000 517.960000 9.655000 519.040000 ;
      RECT 7.060000 513.600000 9.820000 517.960000 ;
      RECT 7.060000 512.520000 9.655000 513.600000 ;
      RECT 7.060000 508.160000 9.820000 512.520000 ;
      RECT 7.060000 507.080000 9.655000 508.160000 ;
      RECT 7.060000 502.720000 9.820000 507.080000 ;
      RECT 7.060000 501.640000 9.655000 502.720000 ;
      RECT 7.060000 497.280000 9.820000 501.640000 ;
      RECT 7.060000 496.200000 9.655000 497.280000 ;
      RECT 7.060000 491.840000 9.820000 496.200000 ;
      RECT 7.060000 490.760000 9.655000 491.840000 ;
      RECT 7.060000 486.400000 9.820000 490.760000 ;
      RECT 7.060000 485.320000 9.655000 486.400000 ;
      RECT 7.060000 480.960000 9.820000 485.320000 ;
      RECT 7.060000 479.880000 9.655000 480.960000 ;
      RECT 7.060000 475.520000 9.820000 479.880000 ;
      RECT 7.060000 474.440000 9.655000 475.520000 ;
      RECT 7.060000 470.080000 9.820000 474.440000 ;
      RECT 7.060000 469.000000 9.655000 470.080000 ;
      RECT 7.060000 464.640000 9.820000 469.000000 ;
      RECT 7.060000 463.560000 9.655000 464.640000 ;
      RECT 7.060000 459.200000 9.820000 463.560000 ;
      RECT 7.060000 458.120000 9.655000 459.200000 ;
      RECT 7.060000 453.760000 9.820000 458.120000 ;
      RECT 7.060000 452.680000 9.655000 453.760000 ;
      RECT 7.060000 448.320000 9.820000 452.680000 ;
      RECT 7.060000 447.240000 9.655000 448.320000 ;
      RECT 7.060000 442.880000 9.820000 447.240000 ;
      RECT 7.060000 441.800000 9.655000 442.880000 ;
      RECT 7.060000 437.440000 9.820000 441.800000 ;
      RECT 7.060000 436.360000 9.655000 437.440000 ;
      RECT 7.060000 432.000000 9.820000 436.360000 ;
      RECT 7.060000 430.920000 9.655000 432.000000 ;
      RECT 7.060000 426.560000 9.820000 430.920000 ;
      RECT 7.060000 425.480000 9.655000 426.560000 ;
      RECT 7.060000 421.120000 9.820000 425.480000 ;
      RECT 7.060000 420.040000 9.655000 421.120000 ;
      RECT 7.060000 415.680000 9.820000 420.040000 ;
      RECT 7.060000 414.600000 9.655000 415.680000 ;
      RECT 7.060000 410.240000 9.820000 414.600000 ;
      RECT 7.060000 409.160000 9.655000 410.240000 ;
      RECT 7.060000 404.800000 9.820000 409.160000 ;
      RECT 7.060000 403.720000 9.655000 404.800000 ;
      RECT 7.060000 399.360000 9.820000 403.720000 ;
      RECT 7.060000 398.280000 9.655000 399.360000 ;
      RECT 7.060000 393.920000 9.820000 398.280000 ;
      RECT 7.060000 392.840000 9.655000 393.920000 ;
      RECT 7.060000 388.480000 9.820000 392.840000 ;
      RECT 7.060000 387.400000 9.655000 388.480000 ;
      RECT 7.060000 383.040000 9.820000 387.400000 ;
      RECT 7.060000 381.960000 9.655000 383.040000 ;
      RECT 7.060000 377.600000 9.820000 381.960000 ;
      RECT 7.060000 376.520000 9.655000 377.600000 ;
      RECT 7.060000 372.160000 9.820000 376.520000 ;
      RECT 7.060000 371.080000 9.655000 372.160000 ;
      RECT 7.060000 366.720000 9.820000 371.080000 ;
      RECT 7.060000 365.640000 9.655000 366.720000 ;
      RECT 7.060000 361.280000 9.820000 365.640000 ;
      RECT 7.060000 360.200000 9.655000 361.280000 ;
      RECT 7.060000 355.840000 9.820000 360.200000 ;
      RECT 7.060000 354.760000 9.655000 355.840000 ;
      RECT 7.060000 350.400000 9.820000 354.760000 ;
      RECT 7.060000 349.320000 9.655000 350.400000 ;
      RECT 7.060000 344.960000 9.820000 349.320000 ;
      RECT 7.060000 343.880000 9.655000 344.960000 ;
      RECT 7.060000 339.520000 9.820000 343.880000 ;
      RECT 7.060000 338.440000 9.655000 339.520000 ;
      RECT 7.060000 334.080000 9.820000 338.440000 ;
      RECT 7.060000 333.000000 9.655000 334.080000 ;
      RECT 7.060000 328.640000 9.820000 333.000000 ;
      RECT 7.060000 327.560000 9.655000 328.640000 ;
      RECT 7.060000 323.200000 9.820000 327.560000 ;
      RECT 7.060000 322.120000 9.655000 323.200000 ;
      RECT 7.060000 317.760000 9.820000 322.120000 ;
      RECT 7.060000 316.680000 9.655000 317.760000 ;
      RECT 7.060000 312.320000 9.820000 316.680000 ;
      RECT 7.060000 311.240000 9.655000 312.320000 ;
      RECT 7.060000 306.880000 9.820000 311.240000 ;
      RECT 7.060000 305.800000 9.655000 306.880000 ;
      RECT 7.060000 301.440000 9.820000 305.800000 ;
      RECT 7.060000 300.360000 9.655000 301.440000 ;
      RECT 7.060000 296.000000 9.820000 300.360000 ;
      RECT 7.060000 294.920000 9.655000 296.000000 ;
      RECT 7.060000 290.560000 9.820000 294.920000 ;
      RECT 7.060000 289.480000 9.655000 290.560000 ;
      RECT 7.060000 285.120000 9.820000 289.480000 ;
      RECT 7.060000 284.040000 9.655000 285.120000 ;
      RECT 7.060000 279.680000 9.820000 284.040000 ;
      RECT 7.060000 278.600000 9.655000 279.680000 ;
      RECT 7.060000 274.240000 9.820000 278.600000 ;
      RECT 7.060000 273.160000 9.655000 274.240000 ;
      RECT 7.060000 268.800000 9.820000 273.160000 ;
      RECT 7.060000 267.720000 9.655000 268.800000 ;
      RECT 7.060000 263.360000 9.820000 267.720000 ;
      RECT 7.060000 262.280000 9.655000 263.360000 ;
      RECT 7.060000 257.920000 9.820000 262.280000 ;
      RECT 7.060000 256.840000 9.655000 257.920000 ;
      RECT 7.060000 252.480000 9.820000 256.840000 ;
      RECT 7.060000 251.400000 9.655000 252.480000 ;
      RECT 7.060000 247.040000 9.820000 251.400000 ;
      RECT 7.060000 245.960000 9.655000 247.040000 ;
      RECT 7.060000 241.600000 9.820000 245.960000 ;
      RECT 7.060000 240.520000 9.655000 241.600000 ;
      RECT 7.060000 236.160000 9.820000 240.520000 ;
      RECT 7.060000 235.080000 9.655000 236.160000 ;
      RECT 7.060000 230.720000 9.820000 235.080000 ;
      RECT 7.060000 229.640000 9.655000 230.720000 ;
      RECT 7.060000 225.280000 9.820000 229.640000 ;
      RECT 7.060000 224.200000 9.655000 225.280000 ;
      RECT 7.060000 219.840000 9.820000 224.200000 ;
      RECT 7.060000 218.760000 9.655000 219.840000 ;
      RECT 7.060000 214.400000 9.820000 218.760000 ;
      RECT 7.060000 213.320000 9.655000 214.400000 ;
      RECT 7.060000 208.960000 9.820000 213.320000 ;
      RECT 7.060000 207.880000 9.655000 208.960000 ;
      RECT 7.060000 203.520000 9.820000 207.880000 ;
      RECT 7.060000 202.440000 9.655000 203.520000 ;
      RECT 7.060000 198.080000 9.820000 202.440000 ;
      RECT 7.060000 197.000000 9.655000 198.080000 ;
      RECT 7.060000 192.640000 9.820000 197.000000 ;
      RECT 7.060000 191.560000 9.655000 192.640000 ;
      RECT 7.060000 187.200000 9.820000 191.560000 ;
      RECT 7.060000 186.120000 9.655000 187.200000 ;
      RECT 7.060000 181.760000 9.820000 186.120000 ;
      RECT 7.060000 180.680000 9.655000 181.760000 ;
      RECT 7.060000 176.320000 9.820000 180.680000 ;
      RECT 7.060000 175.240000 9.655000 176.320000 ;
      RECT 7.060000 170.880000 9.820000 175.240000 ;
      RECT 7.060000 169.800000 9.655000 170.880000 ;
      RECT 7.060000 165.440000 9.820000 169.800000 ;
      RECT 7.060000 164.360000 9.655000 165.440000 ;
      RECT 7.060000 160.000000 9.820000 164.360000 ;
      RECT 7.060000 158.920000 9.655000 160.000000 ;
      RECT 7.060000 154.560000 9.820000 158.920000 ;
      RECT 7.060000 153.480000 9.655000 154.560000 ;
      RECT 7.060000 149.120000 9.820000 153.480000 ;
      RECT 7.060000 148.040000 9.655000 149.120000 ;
      RECT 7.060000 143.680000 9.820000 148.040000 ;
      RECT 7.060000 142.600000 9.655000 143.680000 ;
      RECT 7.060000 138.240000 9.820000 142.600000 ;
      RECT 7.060000 137.160000 9.655000 138.240000 ;
      RECT 7.060000 132.800000 9.820000 137.160000 ;
      RECT 7.060000 131.720000 9.655000 132.800000 ;
      RECT 7.060000 127.360000 9.820000 131.720000 ;
      RECT 7.060000 126.280000 9.655000 127.360000 ;
      RECT 7.060000 121.920000 9.820000 126.280000 ;
      RECT 7.060000 120.840000 9.655000 121.920000 ;
      RECT 7.060000 116.480000 9.820000 120.840000 ;
      RECT 7.060000 115.400000 9.655000 116.480000 ;
      RECT 7.060000 111.040000 9.820000 115.400000 ;
      RECT 7.060000 109.960000 9.655000 111.040000 ;
      RECT 7.060000 105.600000 9.820000 109.960000 ;
      RECT 7.060000 104.520000 9.655000 105.600000 ;
      RECT 7.060000 100.160000 9.820000 104.520000 ;
      RECT 7.060000 99.080000 9.655000 100.160000 ;
      RECT 7.060000 94.720000 9.820000 99.080000 ;
      RECT 7.060000 93.640000 9.655000 94.720000 ;
      RECT 7.060000 89.280000 9.820000 93.640000 ;
      RECT 7.060000 88.200000 9.655000 89.280000 ;
      RECT 7.060000 83.840000 9.820000 88.200000 ;
      RECT 7.060000 82.760000 9.655000 83.840000 ;
      RECT 7.060000 78.400000 9.820000 82.760000 ;
      RECT 7.060000 77.320000 9.655000 78.400000 ;
      RECT 7.060000 72.960000 9.820000 77.320000 ;
      RECT 7.060000 71.880000 9.655000 72.960000 ;
      RECT 7.060000 67.520000 9.820000 71.880000 ;
      RECT 7.060000 66.440000 9.655000 67.520000 ;
      RECT 7.060000 62.080000 9.820000 66.440000 ;
      RECT 7.060000 61.000000 9.655000 62.080000 ;
      RECT 7.060000 56.640000 9.820000 61.000000 ;
      RECT 7.060000 55.560000 9.655000 56.640000 ;
      RECT 7.060000 51.200000 9.820000 55.560000 ;
      RECT 7.060000 50.120000 9.655000 51.200000 ;
      RECT 7.060000 45.760000 9.820000 50.120000 ;
      RECT 7.060000 44.680000 9.655000 45.760000 ;
      RECT 7.060000 40.320000 9.820000 44.680000 ;
      RECT 7.060000 39.240000 9.655000 40.320000 ;
      RECT 7.060000 34.880000 9.820000 39.240000 ;
      RECT 7.060000 33.800000 9.655000 34.880000 ;
      RECT 7.060000 29.440000 9.820000 33.800000 ;
      RECT 7.060000 28.360000 9.655000 29.440000 ;
      RECT 7.060000 24.000000 9.820000 28.360000 ;
      RECT 7.060000 22.920000 9.655000 24.000000 ;
      RECT 7.060000 18.560000 9.820000 22.920000 ;
      RECT 7.060000 17.480000 9.655000 18.560000 ;
      RECT 7.060000 13.120000 9.820000 17.480000 ;
      RECT 7.060000 12.040000 9.655000 13.120000 ;
      RECT 508.620000 5.130000 543.100000 543.460000 ;
      RECT 506.620000 5.130000 506.820000 543.460000 ;
      RECT 463.620000 5.130000 504.820000 543.460000 ;
      RECT 461.620000 5.130000 461.820000 543.460000 ;
      RECT 418.620000 5.130000 459.820000 543.460000 ;
      RECT 416.620000 5.130000 416.820000 543.460000 ;
      RECT 373.620000 5.130000 414.820000 543.460000 ;
      RECT 371.620000 5.130000 371.820000 543.460000 ;
      RECT 328.620000 5.130000 369.820000 543.460000 ;
      RECT 326.620000 5.130000 326.820000 543.460000 ;
      RECT 283.620000 5.130000 324.820000 543.460000 ;
      RECT 281.620000 5.130000 281.820000 543.460000 ;
      RECT 238.620000 5.130000 279.820000 543.460000 ;
      RECT 236.620000 5.130000 236.820000 543.460000 ;
      RECT 193.620000 5.130000 234.820000 543.460000 ;
      RECT 191.620000 5.130000 191.820000 543.460000 ;
      RECT 148.620000 5.130000 189.820000 543.460000 ;
      RECT 146.620000 5.130000 146.820000 543.460000 ;
      RECT 103.620000 5.130000 144.820000 543.460000 ;
      RECT 101.620000 5.130000 101.820000 543.460000 ;
      RECT 58.620000 5.130000 99.820000 543.460000 ;
      RECT 56.620000 5.130000 56.820000 543.460000 ;
      RECT 13.620000 5.130000 54.820000 543.460000 ;
      RECT 11.620000 5.130000 11.820000 543.460000 ;
      RECT 506.620000 2.930000 543.100000 5.130000 ;
      RECT 461.620000 2.930000 504.820000 5.130000 ;
      RECT 416.620000 2.930000 459.820000 5.130000 ;
      RECT 371.620000 2.930000 414.820000 5.130000 ;
      RECT 326.620000 2.930000 369.820000 5.130000 ;
      RECT 281.620000 2.930000 324.820000 5.130000 ;
      RECT 236.620000 2.930000 279.820000 5.130000 ;
      RECT 191.620000 2.930000 234.820000 5.130000 ;
      RECT 146.620000 2.930000 189.820000 5.130000 ;
      RECT 101.620000 2.930000 144.820000 5.130000 ;
      RECT 56.620000 2.930000 99.820000 5.130000 ;
      RECT 11.620000 2.930000 54.820000 5.130000 ;
      RECT 7.060000 2.930000 9.820000 12.040000 ;
      RECT 547.100000 0.000000 550.160000 549.780000 ;
      RECT 544.900000 0.000000 545.300000 549.780000 ;
      RECT 7.060000 0.000000 543.100000 2.930000 ;
      RECT 4.860000 0.000000 5.260000 549.780000 ;
      RECT 0.000000 0.000000 3.060000 549.780000 ;
  END
END flexbex_ibex_core

END LIBRARY
