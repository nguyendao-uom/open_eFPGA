##
## LEF for PtnCells ;
## created by Innovus v19.11-s128_1 on Tue Nov 23 23:09:12 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO S_term_single
  CLASS BLOCK ;
  SIZE 200.100000 BY 30.260000 ;
  FOREIGN S_term_single 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.6048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.696 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 9.240000 29.560000 9.620000 30.260000 ;
    END
  END N1BEG[3]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0871 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.8688 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.104 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 7.860000 29.560000 8.240000 30.260000 ;
    END
  END N1BEG[2]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.061 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 6.480000 29.560000 6.860000 30.260000 ;
    END
  END N1BEG[1]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.313 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 29.560000 5.480000 30.260000 ;
    END
  END N1BEG[0]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1762 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.773 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 21.660000 29.560000 22.040000 30.260000 ;
    END
  END N2BEG[7]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.585 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 19.820000 29.560000 20.200000 30.260000 ;
    END
  END N2BEG[6]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.928 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 18.440000 29.560000 18.820000 30.260000 ;
    END
  END N2BEG[5]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.551 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 17.060000 29.560000 17.440000 30.260000 ;
    END
  END N2BEG[4]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.843 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.107 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 15.680000 29.560000 16.060000 30.260000 ;
    END
  END N2BEG[3]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.251 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 13.840000 29.560000 14.220000 30.260000 ;
    END
  END N2BEG[2]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8222 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.885 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 12.460000 29.560000 12.840000 30.260000 ;
    END
  END N2BEG[1]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4146 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.965 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 11.080000 29.560000 11.460000 30.260000 ;
    END
  END N2BEG[0]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4406 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.977 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 33.620000 29.560000 34.000000 30.260000 ;
    END
  END N2BEGb[7]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0739 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.0768 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.88 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 32.240000 29.560000 32.620000 30.260000 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1764 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.656 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 30.860000 29.560000 31.240000 30.260000 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3362 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 29.020000 29.560000 29.400000 30.260000 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1626 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.705 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 27.640000 29.560000 28.020000 30.260000 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1288 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.418 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 26.260000 29.560000 26.640000 30.260000 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2366 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.957 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 24.420000 29.560000 24.800000 30.260000 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.441 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 23.040000 29.560000 23.420000 30.260000 ;
    END
  END N2BEGb[0]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5358 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.453 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 58.000000 29.560000 58.380000 30.260000 ;
    END
  END N4BEG[15]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6174 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.861 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 56.620000 29.560000 57.000000 30.260000 ;
    END
  END N4BEG[14]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5906 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.845 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 54.780000 29.560000 55.160000 30.260000 ;
    END
  END N4BEG[13]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.551 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 53.400000 29.560000 53.780000 30.260000 ;
    END
  END N4BEG[12]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.77 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.0528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.752 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 52.020000 29.560000 52.400000 30.260000 ;
    END
  END N4BEG[11]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6174 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.861 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 50.180000 29.560000 50.560000 30.260000 ;
    END
  END N4BEG[10]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6526 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.155 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 48.800000 29.560000 49.180000 30.260000 ;
    END
  END N4BEG[9]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.1975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.3738 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.464 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 47.420000 29.560000 47.800000 30.260000 ;
    END
  END N4BEG[8]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2714 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.249 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 45.580000 29.560000 45.960000 30.260000 ;
    END
  END N4BEG[7]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8694 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.121 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 44.200000 29.560000 44.580000 30.260000 ;
    END
  END N4BEG[6]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3458 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.503 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 42.820000 29.560000 43.200000 30.260000 ;
    END
  END N4BEG[5]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.313 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 41.440000 29.560000 41.820000 30.260000 ;
    END
  END N4BEG[4]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2054 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.801 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 39.600000 29.560000 39.980000 30.260000 ;
    END
  END N4BEG[3]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1764 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.656 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 38.220000 29.560000 38.600000 30.260000 ;
    END
  END N4BEG[2]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4077 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.8868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 165.2 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 36.840000 29.560000 37.220000 30.260000 ;
    END
  END N4BEG[1]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.5076 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.648 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 35.000000 29.560000 35.380000 30.260000 ;
    END
  END N4BEG[0]
  PIN NN4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.727 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.409 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 82.380000 29.560000 82.760000 30.260000 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3222 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.503 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 80.540000 29.560000 80.920000 30.260000 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0334 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.059 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 79.160000 29.560000 79.540000 30.260000 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.441 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 77.780000 29.560000 78.160000 30.260000 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.049 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 75.940000 29.560000 76.320000 30.260000 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.848 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 74.560000 29.560000 74.940000 30.260000 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5096 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.322 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 73.180000 29.560000 73.560000 30.260000 ;
    END
  END NN4BEG[9]
  PIN NN4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2655 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.3908 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 103.888 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 71.800000 29.560000 72.180000 30.260000 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5838 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.693 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 69.960000 29.560000 70.340000 30.260000 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8671 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.3316 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.376 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 68.580000 29.560000 68.960000 30.260000 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2865 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.2715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.7368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 116.4 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 67.200000 29.560000 67.580000 30.260000 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.5998 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.773 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 65.360000 29.560000 65.740000 30.260000 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1119 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.4948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.776 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 63.980000 29.560000 64.360000 30.260000 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8385 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.0315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.1938 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 161.504 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 62.600000 29.560000 62.980000 30.260000 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9411 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.6068 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.04 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 60.760000 29.560000 61.140000 30.260000 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.4878 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.213 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 59.380000 29.560000 59.760000 30.260000 ;
    END
  END NN4BEG[0]
  PIN Co
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.928 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 164.260000 29.560000 164.640000 30.260000 ;
    END
  END Co
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.313 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.01939 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.5569 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 88.360000 29.560000 88.740000 30.260000 ;
    END
  END S1END[3]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7703 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.7708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 111.248 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 29.7213 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 157.099 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 86.520000 29.560000 86.900000 30.260000 ;
    END
  END S1END[2]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3838 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.811 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 10.4759 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 50.0047 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 85.140000 29.560000 85.520000 30.260000 ;
    END
  END S1END[1]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.12418 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 9.22626 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 83.760000 29.560000 84.140000 30.260000 ;
    END
  END S1END[0]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5141 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.5018 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.48 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 19.1829 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 101.143 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 112.740000 29.560000 113.120000 30.260000 ;
    END
  END S2MID[7]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0602 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.075 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.02505 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.58519 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 110.900000 29.560000 111.280000 30.260000 ;
    END
  END S2MID[6]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4398 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.973 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.62175 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.9636 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 109.520000 29.560000 109.900000 30.260000 ;
    END
  END S2MID[5]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2827 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.5928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.632 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 16.0378 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 82.3717 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 108.140000 29.560000 108.520000 30.260000 ;
    END
  END S2MID[4]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2941 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.6068 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.04 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 16.962 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 88.7394 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 106.300000 29.560000 106.680000 30.260000 ;
    END
  END S2MID[3]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7586 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.567 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.21589 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.6303 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 104.920000 29.560000 105.300000 30.260000 ;
    END
  END S2MID[2]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.2048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.896 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 29.4827 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 155.203 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 103.540000 29.560000 103.920000 30.260000 ;
    END
  END S2MID[1]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2238 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.011 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 10.9137 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 53.1872 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 101.700000 29.560000 102.080000 30.260000 ;
    END
  END S2MID[0]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0527 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.1025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.1148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 28.2999 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 149.248 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 100.320000 29.560000 100.700000 30.260000 ;
    END
  END S2END[7]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2366 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.957 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.8 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 12.4599 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 98.940000 29.560000 99.320000 30.260000 ;
    END
  END S2END[6]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.313 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.95219 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.31178 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 97.560000 29.560000 97.940000 30.260000 ;
    END
  END S2END[5]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.551 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.0163 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.63232 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 95.720000 29.560000 96.100000 30.260000 ;
    END
  END S2END[4]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3194 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.489 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.13852 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.6155 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 94.340000 29.560000 94.720000 30.260000 ;
    END
  END S2END[3]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.347 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.62721 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 36.7549 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 92.960000 29.560000 93.340000 30.260000 ;
    END
  END S2END[2]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.97024 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.54747 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 91.120000 29.560000 91.500000 30.260000 ;
    END
  END S2END[1]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.835 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.19993 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.3273 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 89.740000 29.560000 90.120000 30.260000 ;
    END
  END S2END[0]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4578 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.063 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.773 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.0337 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 136.660000 29.560000 137.040000 30.260000 ;
    END
  END S4END[15]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.347 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.55515 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 11.3946 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 135.280000 29.560000 135.660000 30.260000 ;
    END
  END S4END[14]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.313 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.95219 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.31178 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 133.900000 29.560000 134.280000 30.260000 ;
    END
  END S4END[13]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7954 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.869 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.11865 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.2121 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 132.060000 29.560000 132.440000 30.260000 ;
    END
  END S4END[12]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.145 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.15663 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.402 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 130.680000 29.560000 131.060000 30.260000 ;
    END
  END S4END[11]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.0376 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 19.8461 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 105.333 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 129.300000 29.560000 129.680000 30.260000 ;
    END
  END S4END[10]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.967 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.0734 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.8269 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 127.460000 29.560000 127.840000 30.260000 ;
    END
  END S4END[9]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.535 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 10.3122 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 50.1798 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 126.080000 29.560000 126.460000 30.260000 ;
    END
  END S4END[8]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.367 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.727 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.43825 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 10.8101 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 124.700000 29.560000 125.080000 30.260000 ;
    END
  END S4END[7]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8906 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.345 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.45306 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.8842 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 123.320000 29.560000 123.700000 30.260000 ;
    END
  END S4END[6]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3194 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.489 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.01764 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.7071 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 121.480000 29.560000 121.860000 30.260000 ;
    END
  END S4END[5]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.88 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.80323 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.635 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 120.100000 29.560000 120.480000 30.260000 ;
    END
  END S4END[4]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.115 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.467 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.0699 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.9684 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 118.720000 29.560000 119.100000 30.260000 ;
    END
  END S4END[3]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5834 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.691 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.22687 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.5865 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 116.880000 29.560000 117.260000 30.260000 ;
    END
  END S4END[2]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.479 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.287 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.41347 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.6862 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 115.500000 29.560000 115.880000 30.260000 ;
    END
  END S4END[1]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.917 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.359 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.43919 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.6559 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 114.120000 29.560000 114.500000 30.260000 ;
    END
  END S4END[0]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.967 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.74465 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.1832 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 161.040000 29.560000 161.420000 30.260000 ;
    END
  END SS4END[15]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8218 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.883 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.9138 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.1199 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 159.660000 29.560000 160.040000 30.260000 ;
    END
  END SS4END[14]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.823 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.46276 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 10.9327 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 157.820000 29.560000 158.200000 30.260000 ;
    END
  END SS4END[13]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.313 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.45306 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 10.7253 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 156.440000 29.560000 156.820000 30.260000 ;
    END
  END SS4END[12]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2974 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.261 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.98936 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.1037 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 155.060000 29.560000 155.440000 30.260000 ;
    END
  END SS4END[11]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.251 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.55024 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.0788 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 153.680000 29.560000 154.060000 30.260000 ;
    END
  END SS4END[10]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1725 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.7648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.216 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 13.4743 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 70.4741 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 151.840000 29.560000 152.220000 30.260000 ;
    END
  END SS4END[9]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7703 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.3688 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.104 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 24.8228 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 131.079 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 150.460000 29.560000 150.840000 30.260000 ;
    END
  END SS4END[8]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.347 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.03475 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.79259 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 149.080000 29.560000 149.460000 30.260000 ;
    END
  END SS4END[7]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5168 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.476 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.03993 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.8249 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 147.240000 29.560000 147.620000 30.260000 ;
    END
  END SS4END[6]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7742 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.645 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.83138 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.6168 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 145.860000 29.560000 146.240000 30.260000 ;
    END
  END SS4END[5]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.305 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.417 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.43542 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 45.796 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 144.480000 29.560000 144.860000 30.260000 ;
    END
  END SS4END[4]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.428 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.39616 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.6061 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 142.640000 29.560000 143.020000 30.260000 ;
    END
  END SS4END[3]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.025 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.73145 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.1172 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 141.260000 29.560000 141.640000 30.260000 ;
    END
  END SS4END[2]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0736 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.25 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.06007 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.90572 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 139.880000 29.560000 140.260000 30.260000 ;
    END
  END SS4END[1]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0814 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.299 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.24525 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.8451 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 138.500000 29.560000 138.880000 30.260000 ;
    END
  END SS4END[0]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.152 LAYER met3  ;
    ANTENNAMAXAREACAR 2.16855 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 9.50868 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.0793403 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 0.000000 5.480000 0.700000 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1552 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.766 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 162.420000 29.560000 162.800000 30.260000 ;
    END
  END UserCLKo
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3666 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.725 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.47838 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.0108 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 194.620000 0.000000 195.000000 0.700000 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0974 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.379 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.94552 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 27.0552 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 184.960000 0.000000 185.340000 0.700000 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6522 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.153 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.22216 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 28.736 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 175.300000 0.000000 175.680000 0.700000 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.257 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.177 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.35104 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.6781 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 166.100000 0.000000 166.480000 0.700000 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.068 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.45852 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.2155 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 156.440000 0.000000 156.820000 0.700000 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.781 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.797 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.50707 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.1542 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 147.240000 0.000000 147.620000 0.700000 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0839 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.5028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.152 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 14.3615 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 75.332 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 137.580000 0.000000 137.960000 0.700000 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.869 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.119 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.32417 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.1717 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 127.920000 0.000000 128.300000 0.700000 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.082 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.1132 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.8256 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 118.720000 0.000000 119.100000 0.700000 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3444 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.604 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.96444 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.5185 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 109.060000 0.000000 109.440000 0.700000 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.976 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.47758 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.9387 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 99.400000 0.000000 99.780000 0.700000 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9088 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.308 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.37778 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.4263 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 90.200000 0.000000 90.580000 0.700000 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.525 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.65724 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.7461 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 80.540000 0.000000 80.920000 0.700000 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5834 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.691 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.93953 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.2485 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 71.340000 0.000000 71.720000 0.700000 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6646 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.097 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.93818 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.1508 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 61.680000 0.000000 62.060000 0.700000 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9317 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.5448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.376 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 36.0007 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 189.883 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 52.480000 0.000000 52.860000 0.700000 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2362 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.955 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.47192 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.9104 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 42.820000 0.000000 43.200000 0.700000 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5358 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.453 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.87542 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.9279 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 33.160000 0.000000 33.540000 0.700000 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9017 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.1098 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.056 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 22.0978 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 116.531 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 23.960000 0.000000 24.340000 0.700000 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5972 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.868 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.08828 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.7556 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 14.300000 0.000000 14.680000 0.700000 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6526 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.155 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 194.160000 29.560000 194.540000 30.260000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.585 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 192.780000 29.560000 193.160000 30.260000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.367 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.727 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 191.400000 29.560000 191.780000 30.260000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.061 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 190.020000 29.560000 190.400000 30.260000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8122 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.953 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 188.180000 29.560000 188.560000 30.260000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4314 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.049 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 186.800000 29.560000 187.180000 30.260000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5362 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.455 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 185.420000 29.560000 185.800000 30.260000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5362 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.455 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 183.580000 29.560000 183.960000 30.260000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6526 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.155 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 182.200000 29.560000 182.580000 30.260000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.585 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 180.820000 29.560000 181.200000 30.260000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4266 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.907 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 179.440000 29.560000 179.820000 30.260000 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5362 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.455 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 177.600000 29.560000 177.980000 30.260000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.154 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 176.220000 29.560000 176.600000 30.260000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.548 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 174.840000 29.560000 175.220000 30.260000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6856 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.202 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 173.000000 29.560000 173.380000 30.260000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7455 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.2688 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.904 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 171.620000 29.560000 172.000000 30.260000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2714 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.249 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 170.240000 29.560000 170.620000 30.260000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3433 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5555 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.7308 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 168.400000 29.560000 168.780000 30.260000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.205 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 167.020000 29.560000 167.400000 30.260000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6214 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.999 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 165.640000 29.560000 166.020000 30.260000 ;
    END
  END FrameStrobe_O[0]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 198.900000 25.700000 200.100000 26.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 25.700000 1.200000 26.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.900000 2.850000 200.100000 4.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 1.200000 4.050000 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.070000 29.060000 197.270000 30.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.070000 0.000000 197.270000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 29.060000 4.030000 30.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 0.000000 4.030000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 200.100000 4.050000 ;
        RECT 0.000000 25.700000 200.100000 26.900000 ;
        RECT 7.060000 4.860000 8.260000 5.340000 ;
        RECT 2.830000 4.860000 4.030000 5.340000 ;
        RECT 7.060000 10.300000 8.260000 10.780000 ;
        RECT 2.830000 10.300000 4.030000 10.780000 ;
        RECT 52.060000 10.300000 53.260000 10.780000 ;
        RECT 97.060000 10.300000 98.260000 10.780000 ;
        RECT 97.060000 4.860000 98.260000 5.340000 ;
        RECT 52.060000 4.860000 53.260000 5.340000 ;
        RECT 142.060000 10.300000 143.260000 10.780000 ;
        RECT 142.060000 4.860000 143.260000 5.340000 ;
        RECT 187.060000 4.860000 188.260000 5.340000 ;
        RECT 187.060000 10.300000 188.260000 10.780000 ;
        RECT 196.070000 10.300000 197.270000 10.780000 ;
        RECT 196.070000 4.860000 197.270000 5.340000 ;
        RECT 2.830000 21.180000 4.030000 21.660000 ;
        RECT 7.060000 21.180000 8.260000 21.660000 ;
        RECT 7.060000 15.740000 8.260000 16.220000 ;
        RECT 2.830000 15.740000 4.030000 16.220000 ;
        RECT 52.060000 21.180000 53.260000 21.660000 ;
        RECT 97.060000 21.180000 98.260000 21.660000 ;
        RECT 97.060000 15.740000 98.260000 16.220000 ;
        RECT 52.060000 15.740000 53.260000 16.220000 ;
        RECT 142.060000 21.180000 143.260000 21.660000 ;
        RECT 142.060000 15.740000 143.260000 16.220000 ;
        RECT 187.060000 15.740000 188.260000 16.220000 ;
        RECT 187.060000 21.180000 188.260000 21.660000 ;
        RECT 196.070000 21.180000 197.270000 21.660000 ;
        RECT 196.070000 15.740000 197.270000 16.220000 ;
      LAYER met4 ;
        RECT 187.060000 2.850000 188.260000 26.900000 ;
        RECT 142.060000 2.850000 143.260000 26.900000 ;
        RECT 97.060000 2.850000 98.260000 26.900000 ;
        RECT 52.060000 2.850000 53.260000 26.900000 ;
        RECT 7.060000 2.850000 8.260000 26.900000 ;
        RECT 196.070000 0.000000 197.270000 30.260000 ;
        RECT 2.830000 0.000000 4.030000 30.260000 ;
    END
# end of P/G power stripe data as pin

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 198.900000 27.500000 200.100000 28.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 27.500000 1.200000 28.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.900000 1.050000 200.100000 2.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 1.200000 2.250000 ;
    END
    PORT
      LAYER met4 ;
        RECT 197.870000 29.060000 199.070000 30.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 197.870000 0.000000 199.070000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 29.060000 2.230000 30.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 0.000000 2.230000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 200.100000 2.250000 ;
        RECT 0.000000 27.500000 200.100000 28.700000 ;
        RECT 1.030000 7.580000 2.230000 8.060000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 1.030000 13.020000 2.230000 13.500000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 50.060000 13.020000 51.260000 13.500000 ;
        RECT 95.060000 13.020000 96.260000 13.500000 ;
        RECT 50.060000 7.580000 51.260000 8.060000 ;
        RECT 95.060000 7.580000 96.260000 8.060000 ;
        RECT 140.060000 13.020000 141.260000 13.500000 ;
        RECT 140.060000 7.580000 141.260000 8.060000 ;
        RECT 185.060000 7.580000 186.260000 8.060000 ;
        RECT 185.060000 13.020000 186.260000 13.500000 ;
        RECT 197.870000 7.580000 199.070000 8.060000 ;
        RECT 197.870000 13.020000 199.070000 13.500000 ;
        RECT 1.030000 18.460000 2.230000 18.940000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 1.030000 23.900000 2.230000 24.380000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
        RECT 50.060000 23.900000 51.260000 24.380000 ;
        RECT 95.060000 23.900000 96.260000 24.380000 ;
        RECT 50.060000 18.460000 51.260000 18.940000 ;
        RECT 95.060000 18.460000 96.260000 18.940000 ;
        RECT 140.060000 23.900000 141.260000 24.380000 ;
        RECT 140.060000 18.460000 141.260000 18.940000 ;
        RECT 185.060000 18.460000 186.260000 18.940000 ;
        RECT 185.060000 23.900000 186.260000 24.380000 ;
        RECT 197.870000 18.460000 199.070000 18.940000 ;
        RECT 197.870000 23.900000 199.070000 24.380000 ;
      LAYER met4 ;
        RECT 185.060000 1.050000 186.260000 28.700000 ;
        RECT 140.060000 1.050000 141.260000 28.700000 ;
        RECT 95.060000 1.050000 96.260000 28.700000 ;
        RECT 50.060000 1.050000 51.260000 28.700000 ;
        RECT 5.060000 1.050000 6.260000 28.700000 ;
        RECT 197.870000 0.000000 199.070000 30.260000 ;
        RECT 1.030000 0.000000 2.230000 30.260000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
    END
# end of P/G power stripe data as pin

  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 200.100000 30.260000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 200.100000 30.260000 ;
    LAYER met2 ;
      RECT 194.680000 29.420000 200.100000 30.260000 ;
      RECT 193.300000 29.420000 194.020000 30.260000 ;
      RECT 191.920000 29.420000 192.640000 30.260000 ;
      RECT 190.540000 29.420000 191.260000 30.260000 ;
      RECT 188.700000 29.420000 189.880000 30.260000 ;
      RECT 187.320000 29.420000 188.040000 30.260000 ;
      RECT 185.940000 29.420000 186.660000 30.260000 ;
      RECT 184.100000 29.420000 185.280000 30.260000 ;
      RECT 182.720000 29.420000 183.440000 30.260000 ;
      RECT 181.340000 29.420000 182.060000 30.260000 ;
      RECT 179.960000 29.420000 180.680000 30.260000 ;
      RECT 178.120000 29.420000 179.300000 30.260000 ;
      RECT 176.740000 29.420000 177.460000 30.260000 ;
      RECT 175.360000 29.420000 176.080000 30.260000 ;
      RECT 173.520000 29.420000 174.700000 30.260000 ;
      RECT 172.140000 29.420000 172.860000 30.260000 ;
      RECT 170.760000 29.420000 171.480000 30.260000 ;
      RECT 168.920000 29.420000 170.100000 30.260000 ;
      RECT 167.540000 29.420000 168.260000 30.260000 ;
      RECT 166.160000 29.420000 166.880000 30.260000 ;
      RECT 164.780000 29.420000 165.500000 30.260000 ;
      RECT 162.940000 29.420000 164.120000 30.260000 ;
      RECT 161.560000 29.420000 162.280000 30.260000 ;
      RECT 160.180000 29.420000 160.900000 30.260000 ;
      RECT 158.340000 29.420000 159.520000 30.260000 ;
      RECT 156.960000 29.420000 157.680000 30.260000 ;
      RECT 155.580000 29.420000 156.300000 30.260000 ;
      RECT 154.200000 29.420000 154.920000 30.260000 ;
      RECT 152.360000 29.420000 153.540000 30.260000 ;
      RECT 150.980000 29.420000 151.700000 30.260000 ;
      RECT 149.600000 29.420000 150.320000 30.260000 ;
      RECT 147.760000 29.420000 148.940000 30.260000 ;
      RECT 146.380000 29.420000 147.100000 30.260000 ;
      RECT 145.000000 29.420000 145.720000 30.260000 ;
      RECT 143.160000 29.420000 144.340000 30.260000 ;
      RECT 141.780000 29.420000 142.500000 30.260000 ;
      RECT 140.400000 29.420000 141.120000 30.260000 ;
      RECT 139.020000 29.420000 139.740000 30.260000 ;
      RECT 137.180000 29.420000 138.360000 30.260000 ;
      RECT 135.800000 29.420000 136.520000 30.260000 ;
      RECT 134.420000 29.420000 135.140000 30.260000 ;
      RECT 132.580000 29.420000 133.760000 30.260000 ;
      RECT 131.200000 29.420000 131.920000 30.260000 ;
      RECT 129.820000 29.420000 130.540000 30.260000 ;
      RECT 127.980000 29.420000 129.160000 30.260000 ;
      RECT 126.600000 29.420000 127.320000 30.260000 ;
      RECT 125.220000 29.420000 125.940000 30.260000 ;
      RECT 123.840000 29.420000 124.560000 30.260000 ;
      RECT 122.000000 29.420000 123.180000 30.260000 ;
      RECT 120.620000 29.420000 121.340000 30.260000 ;
      RECT 119.240000 29.420000 119.960000 30.260000 ;
      RECT 117.400000 29.420000 118.580000 30.260000 ;
      RECT 116.020000 29.420000 116.740000 30.260000 ;
      RECT 114.640000 29.420000 115.360000 30.260000 ;
      RECT 113.260000 29.420000 113.980000 30.260000 ;
      RECT 111.420000 29.420000 112.600000 30.260000 ;
      RECT 110.040000 29.420000 110.760000 30.260000 ;
      RECT 108.660000 29.420000 109.380000 30.260000 ;
      RECT 106.820000 29.420000 108.000000 30.260000 ;
      RECT 105.440000 29.420000 106.160000 30.260000 ;
      RECT 104.060000 29.420000 104.780000 30.260000 ;
      RECT 102.220000 29.420000 103.400000 30.260000 ;
      RECT 100.840000 29.420000 101.560000 30.260000 ;
      RECT 99.460000 29.420000 100.180000 30.260000 ;
      RECT 98.080000 29.420000 98.800000 30.260000 ;
      RECT 96.240000 29.420000 97.420000 30.260000 ;
      RECT 94.860000 29.420000 95.580000 30.260000 ;
      RECT 93.480000 29.420000 94.200000 30.260000 ;
      RECT 91.640000 29.420000 92.820000 30.260000 ;
      RECT 90.260000 29.420000 90.980000 30.260000 ;
      RECT 88.880000 29.420000 89.600000 30.260000 ;
      RECT 87.040000 29.420000 88.220000 30.260000 ;
      RECT 85.660000 29.420000 86.380000 30.260000 ;
      RECT 84.280000 29.420000 85.000000 30.260000 ;
      RECT 82.900000 29.420000 83.620000 30.260000 ;
      RECT 81.060000 29.420000 82.240000 30.260000 ;
      RECT 79.680000 29.420000 80.400000 30.260000 ;
      RECT 78.300000 29.420000 79.020000 30.260000 ;
      RECT 76.460000 29.420000 77.640000 30.260000 ;
      RECT 75.080000 29.420000 75.800000 30.260000 ;
      RECT 73.700000 29.420000 74.420000 30.260000 ;
      RECT 72.320000 29.420000 73.040000 30.260000 ;
      RECT 70.480000 29.420000 71.660000 30.260000 ;
      RECT 69.100000 29.420000 69.820000 30.260000 ;
      RECT 67.720000 29.420000 68.440000 30.260000 ;
      RECT 65.880000 29.420000 67.060000 30.260000 ;
      RECT 64.500000 29.420000 65.220000 30.260000 ;
      RECT 63.120000 29.420000 63.840000 30.260000 ;
      RECT 61.280000 29.420000 62.460000 30.260000 ;
      RECT 59.900000 29.420000 60.620000 30.260000 ;
      RECT 58.520000 29.420000 59.240000 30.260000 ;
      RECT 57.140000 29.420000 57.860000 30.260000 ;
      RECT 55.300000 29.420000 56.480000 30.260000 ;
      RECT 53.920000 29.420000 54.640000 30.260000 ;
      RECT 52.540000 29.420000 53.260000 30.260000 ;
      RECT 50.700000 29.420000 51.880000 30.260000 ;
      RECT 49.320000 29.420000 50.040000 30.260000 ;
      RECT 47.940000 29.420000 48.660000 30.260000 ;
      RECT 46.100000 29.420000 47.280000 30.260000 ;
      RECT 44.720000 29.420000 45.440000 30.260000 ;
      RECT 43.340000 29.420000 44.060000 30.260000 ;
      RECT 41.960000 29.420000 42.680000 30.260000 ;
      RECT 40.120000 29.420000 41.300000 30.260000 ;
      RECT 38.740000 29.420000 39.460000 30.260000 ;
      RECT 37.360000 29.420000 38.080000 30.260000 ;
      RECT 35.520000 29.420000 36.700000 30.260000 ;
      RECT 34.140000 29.420000 34.860000 30.260000 ;
      RECT 32.760000 29.420000 33.480000 30.260000 ;
      RECT 31.380000 29.420000 32.100000 30.260000 ;
      RECT 29.540000 29.420000 30.720000 30.260000 ;
      RECT 28.160000 29.420000 28.880000 30.260000 ;
      RECT 26.780000 29.420000 27.500000 30.260000 ;
      RECT 24.940000 29.420000 26.120000 30.260000 ;
      RECT 23.560000 29.420000 24.280000 30.260000 ;
      RECT 22.180000 29.420000 22.900000 30.260000 ;
      RECT 20.340000 29.420000 21.520000 30.260000 ;
      RECT 18.960000 29.420000 19.680000 30.260000 ;
      RECT 17.580000 29.420000 18.300000 30.260000 ;
      RECT 16.200000 29.420000 16.920000 30.260000 ;
      RECT 14.360000 29.420000 15.540000 30.260000 ;
      RECT 12.980000 29.420000 13.700000 30.260000 ;
      RECT 11.600000 29.420000 12.320000 30.260000 ;
      RECT 9.760000 29.420000 10.940000 30.260000 ;
      RECT 8.380000 29.420000 9.100000 30.260000 ;
      RECT 7.000000 29.420000 7.720000 30.260000 ;
      RECT 5.620000 29.420000 6.340000 30.260000 ;
      RECT 0.000000 29.420000 4.960000 30.260000 ;
      RECT 0.000000 0.840000 200.100000 29.420000 ;
      RECT 195.140000 0.000000 200.100000 0.840000 ;
      RECT 185.480000 0.000000 194.480000 0.840000 ;
      RECT 175.820000 0.000000 184.820000 0.840000 ;
      RECT 166.620000 0.000000 175.160000 0.840000 ;
      RECT 156.960000 0.000000 165.960000 0.840000 ;
      RECT 147.760000 0.000000 156.300000 0.840000 ;
      RECT 138.100000 0.000000 147.100000 0.840000 ;
      RECT 128.440000 0.000000 137.440000 0.840000 ;
      RECT 119.240000 0.000000 127.780000 0.840000 ;
      RECT 109.580000 0.000000 118.580000 0.840000 ;
      RECT 99.920000 0.000000 108.920000 0.840000 ;
      RECT 90.720000 0.000000 99.260000 0.840000 ;
      RECT 81.060000 0.000000 90.060000 0.840000 ;
      RECT 71.860000 0.000000 80.400000 0.840000 ;
      RECT 62.200000 0.000000 71.200000 0.840000 ;
      RECT 53.000000 0.000000 61.540000 0.840000 ;
      RECT 43.340000 0.000000 52.340000 0.840000 ;
      RECT 33.680000 0.000000 42.680000 0.840000 ;
      RECT 24.480000 0.000000 33.020000 0.840000 ;
      RECT 14.820000 0.000000 23.820000 0.840000 ;
      RECT 5.620000 0.000000 14.160000 0.840000 ;
      RECT 0.000000 0.000000 4.960000 0.840000 ;
    LAYER met3 ;
      RECT 0.000000 29.000000 200.100000 30.260000 ;
      RECT 0.000000 24.680000 200.100000 25.400000 ;
      RECT 199.370000 23.600000 200.100000 24.680000 ;
      RECT 186.560000 23.600000 197.570000 24.680000 ;
      RECT 141.560000 23.600000 184.760000 24.680000 ;
      RECT 96.560000 23.600000 139.760000 24.680000 ;
      RECT 51.560000 23.600000 94.760000 24.680000 ;
      RECT 6.560000 23.600000 49.760000 24.680000 ;
      RECT 2.530000 23.600000 4.595000 24.680000 ;
      RECT 0.000000 23.600000 0.730000 24.680000 ;
      RECT 0.000000 21.960000 200.100000 23.600000 ;
      RECT 197.570000 20.880000 200.100000 21.960000 ;
      RECT 188.560000 20.880000 195.770000 21.960000 ;
      RECT 143.560000 20.880000 186.760000 21.960000 ;
      RECT 98.560000 20.880000 141.760000 21.960000 ;
      RECT 53.560000 20.880000 96.760000 21.960000 ;
      RECT 8.560000 20.880000 51.760000 21.960000 ;
      RECT 4.330000 20.880000 6.760000 21.960000 ;
      RECT 0.000000 20.880000 2.530000 21.960000 ;
      RECT 0.000000 19.240000 200.100000 20.880000 ;
      RECT 199.370000 18.160000 200.100000 19.240000 ;
      RECT 186.560000 18.160000 197.570000 19.240000 ;
      RECT 141.560000 18.160000 184.760000 19.240000 ;
      RECT 96.560000 18.160000 139.760000 19.240000 ;
      RECT 51.560000 18.160000 94.760000 19.240000 ;
      RECT 6.560000 18.160000 49.760000 19.240000 ;
      RECT 2.530000 18.160000 4.595000 19.240000 ;
      RECT 0.000000 18.160000 0.730000 19.240000 ;
      RECT 0.000000 16.520000 200.100000 18.160000 ;
      RECT 197.570000 15.440000 200.100000 16.520000 ;
      RECT 188.560000 15.440000 195.770000 16.520000 ;
      RECT 143.560000 15.440000 186.760000 16.520000 ;
      RECT 98.560000 15.440000 141.760000 16.520000 ;
      RECT 53.560000 15.440000 96.760000 16.520000 ;
      RECT 8.560000 15.440000 51.760000 16.520000 ;
      RECT 4.330000 15.440000 6.760000 16.520000 ;
      RECT 0.000000 15.440000 2.530000 16.520000 ;
      RECT 0.000000 13.800000 200.100000 15.440000 ;
      RECT 199.370000 12.720000 200.100000 13.800000 ;
      RECT 186.560000 12.720000 197.570000 13.800000 ;
      RECT 141.560000 12.720000 184.760000 13.800000 ;
      RECT 96.560000 12.720000 139.760000 13.800000 ;
      RECT 51.560000 12.720000 94.760000 13.800000 ;
      RECT 6.560000 12.720000 49.760000 13.800000 ;
      RECT 2.530000 12.720000 4.595000 13.800000 ;
      RECT 0.000000 12.720000 0.730000 13.800000 ;
      RECT 0.000000 11.080000 200.100000 12.720000 ;
      RECT 197.570000 10.000000 200.100000 11.080000 ;
      RECT 188.560000 10.000000 195.770000 11.080000 ;
      RECT 143.560000 10.000000 186.760000 11.080000 ;
      RECT 98.560000 10.000000 141.760000 11.080000 ;
      RECT 53.560000 10.000000 96.760000 11.080000 ;
      RECT 8.560000 10.000000 51.760000 11.080000 ;
      RECT 4.330000 10.000000 6.760000 11.080000 ;
      RECT 0.000000 10.000000 2.530000 11.080000 ;
      RECT 0.000000 8.360000 200.100000 10.000000 ;
      RECT 199.370000 7.280000 200.100000 8.360000 ;
      RECT 186.560000 7.280000 197.570000 8.360000 ;
      RECT 141.560000 7.280000 184.760000 8.360000 ;
      RECT 96.560000 7.280000 139.760000 8.360000 ;
      RECT 51.560000 7.280000 94.760000 8.360000 ;
      RECT 6.560000 7.280000 49.760000 8.360000 ;
      RECT 2.530000 7.280000 4.595000 8.360000 ;
      RECT 0.000000 7.280000 0.730000 8.360000 ;
      RECT 0.000000 5.640000 200.100000 7.280000 ;
      RECT 197.570000 4.560000 200.100000 5.640000 ;
      RECT 188.560000 4.560000 195.770000 5.640000 ;
      RECT 143.560000 4.560000 186.760000 5.640000 ;
      RECT 98.560000 4.560000 141.760000 5.640000 ;
      RECT 53.560000 4.560000 96.760000 5.640000 ;
      RECT 8.560000 4.560000 51.760000 5.640000 ;
      RECT 4.330000 4.560000 6.760000 5.640000 ;
      RECT 0.000000 4.560000 2.530000 5.640000 ;
      RECT 0.000000 4.350000 200.100000 4.560000 ;
      RECT 0.000000 0.000000 200.100000 0.750000 ;
    LAYER met4 ;
      RECT 4.330000 29.000000 195.770000 30.260000 ;
      RECT 186.560000 27.200000 195.770000 29.000000 ;
      RECT 141.560000 27.200000 184.760000 29.000000 ;
      RECT 96.560000 27.200000 139.760000 29.000000 ;
      RECT 51.560000 27.200000 94.760000 29.000000 ;
      RECT 6.560000 27.200000 49.760000 29.000000 ;
      RECT 4.330000 24.680000 4.760000 29.000000 ;
      RECT 4.330000 23.600000 4.595000 24.680000 ;
      RECT 4.330000 19.240000 4.760000 23.600000 ;
      RECT 4.330000 18.160000 4.595000 19.240000 ;
      RECT 4.330000 13.800000 4.760000 18.160000 ;
      RECT 4.330000 12.720000 4.595000 13.800000 ;
      RECT 4.330000 8.360000 4.760000 12.720000 ;
      RECT 4.330000 7.280000 4.595000 8.360000 ;
      RECT 188.560000 2.550000 195.770000 27.200000 ;
      RECT 186.560000 2.550000 186.760000 27.200000 ;
      RECT 143.560000 2.550000 184.760000 27.200000 ;
      RECT 141.560000 2.550000 141.760000 27.200000 ;
      RECT 98.560000 2.550000 139.760000 27.200000 ;
      RECT 96.560000 2.550000 96.760000 27.200000 ;
      RECT 53.560000 2.550000 94.760000 27.200000 ;
      RECT 51.560000 2.550000 51.760000 27.200000 ;
      RECT 8.560000 2.550000 49.760000 27.200000 ;
      RECT 6.560000 2.550000 6.760000 27.200000 ;
      RECT 186.560000 0.750000 195.770000 2.550000 ;
      RECT 141.560000 0.750000 184.760000 2.550000 ;
      RECT 96.560000 0.750000 139.760000 2.550000 ;
      RECT 51.560000 0.750000 94.760000 2.550000 ;
      RECT 6.560000 0.750000 49.760000 2.550000 ;
      RECT 4.330000 0.750000 4.760000 7.280000 ;
      RECT 199.370000 0.000000 200.100000 30.260000 ;
      RECT 4.330000 0.000000 195.770000 0.750000 ;
      RECT 0.000000 0.000000 0.730000 30.260000 ;
  END
END S_term_single

END LIBRARY
