##
## LEF for PtnCells ;
## created by Innovus v19.11-s128_1 on Thu Dec  2 18:40:22 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO W_CPU_IO
  CLASS BLOCK ;
  SIZE 40.020000 BY 200.260000 ;
  FOREIGN W_CPU_IO 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1766 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.3468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.32 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 80.720000 40.020000 81.100000 ;
    END
  END E1BEG[3]
  PIN E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2576 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.0768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 96.88 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 79.500000 40.020000 79.880000 ;
    END
  END E1BEG[2]
  PIN E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 77.670000 40.020000 78.050000 ;
    END
  END E1BEG[1]
  PIN E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.9204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.904 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 76.450000 40.020000 76.830000 ;
    END
  END E1BEG[0]
  PIN E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 92.920000 40.020000 93.300000 ;
    END
  END E2BEG[7]
  PIN E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8216 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.04 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.0768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 96.88 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 91.090000 40.020000 91.470000 ;
    END
  END E2BEG[6]
  PIN E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 89.870000 40.020000 90.250000 ;
    END
  END E2BEG[5]
  PIN E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.712 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 88.040000 40.020000 88.420000 ;
    END
  END E2BEG[4]
  PIN E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 86.820000 40.020000 87.200000 ;
    END
  END E2BEG[3]
  PIN E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.3874 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.728 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 84.990000 40.020000 85.370000 ;
    END
  END E2BEG[2]
  PIN E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 83.770000 40.020000 84.150000 ;
    END
  END E2BEG[1]
  PIN E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 81.940000 40.020000 82.320000 ;
    END
  END E2BEG[0]
  PIN E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 104.510000 40.020000 104.890000 ;
    END
  END E2BEGb[7]
  PIN E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0156 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.9308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 106.768 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 103.290000 40.020000 103.670000 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0376 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.9548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 90.896 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 101.460000 40.020000 101.840000 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 100.240000 40.020000 100.620000 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 98.410000 40.020000 98.790000 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.392 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.1618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 92 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 97.190000 40.020000 97.570000 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 95.360000 40.020000 95.740000 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 94.140000 40.020000 94.520000 ;
    END
  END E2BEGb[0]
  PIN EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 128.300000 40.020000 128.680000 ;
    END
  END EE4BEG[15]
  PIN EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5396 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.1768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 124.08 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 127.080000 40.020000 127.460000 ;
    END
  END EE4BEG[14]
  PIN EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 125.250000 40.020000 125.630000 ;
    END
  END EE4BEG[13]
  PIN EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1134 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.4 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.0658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 107.488 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 124.030000 40.020000 124.410000 ;
    END
  END EE4BEG[12]
  PIN EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8514 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.536 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 122.200000 40.020000 122.580000 ;
    END
  END EE4BEG[11]
  PIN EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0636 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.664 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.6018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.68 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 120.980000 40.020000 121.360000 ;
    END
  END EE4BEG[10]
  PIN EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 119.150000 40.020000 119.530000 ;
    END
  END EE4BEG[9]
  PIN EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3726 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.9158 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 58.688 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 117.930000 40.020000 118.310000 ;
    END
  END EE4BEG[8]
  PIN EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.2468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 87.12 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 116.710000 40.020000 117.090000 ;
    END
  END EE4BEG[7]
  PIN EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 114.880000 40.020000 115.260000 ;
    END
  END EE4BEG[6]
  PIN EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 113.660000 40.020000 114.040000 ;
    END
  END EE4BEG[5]
  PIN EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 111.830000 40.020000 112.210000 ;
    END
  END EE4BEG[4]
  PIN EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 110.610000 40.020000 110.990000 ;
    END
  END EE4BEG[3]
  PIN EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 108.780000 40.020000 109.160000 ;
    END
  END EE4BEG[2]
  PIN EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.8164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.016 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 107.560000 40.020000 107.940000 ;
    END
  END EE4BEG[1]
  PIN EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 105.730000 40.020000 106.110000 ;
    END
  END EE4BEG[0]
  PIN E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 145.990000 40.020000 146.370000 ;
    END
  END E6BEG[11]
  PIN E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.656 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 144.770000 40.020000 145.150000 ;
    END
  END E6BEG[10]
  PIN E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3354 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.784 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 143.550000 40.020000 143.930000 ;
    END
  END E6BEG[9]
  PIN E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2006 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.4738 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.664 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 141.720000 40.020000 142.100000 ;
    END
  END E6BEG[8]
  PIN E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 140.500000 40.020000 140.880000 ;
    END
  END E6BEG[7]
  PIN E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3174 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 138.670000 40.020000 139.050000 ;
    END
  END E6BEG[6]
  PIN E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 137.450000 40.020000 137.830000 ;
    END
  END E6BEG[5]
  PIN E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 135.620000 40.020000 136.000000 ;
    END
  END E6BEG[4]
  PIN E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 134.400000 40.020000 134.780000 ;
    END
  END E6BEG[3]
  PIN E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.539 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.3428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 71.632 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 132.570000 40.020000 132.950000 ;
    END
  END E6BEG[2]
  PIN E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 131.350000 40.020000 131.730000 ;
    END
  END E6BEG[1]
  PIN E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 130.130000 40.020000 130.510000 ;
    END
  END E6BEG[0]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 7.09751 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 34.2882 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 9.350000 40.020000 9.730000 ;
    END
  END W1END[3]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 4.70976 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 22.0148 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 7.520000 40.020000 7.900000 ;
    END
  END W1END[2]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.656 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 6.47609 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 31.5529 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 6.300000 40.020000 6.680000 ;
    END
  END W1END[1]
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 2.6598 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 12.0377 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 5.080000 40.020000 5.460000 ;
    END
  END W1END[0]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 39.320000 20.940000 40.020000 21.320000 ;
    END
  END W2MID[7]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 7.31488 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 35.6229 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 19.720000 40.020000 20.100000 ;
    END
  END W2MID[6]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 4.63771 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 21.7226 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 17.890000 40.020000 18.270000 ;
    END
  END W2MID[5]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 39.320000 16.670000 40.020000 17.050000 ;
    END
  END W2MID[4]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 39.320000 15.450000 40.020000 15.830000 ;
    END
  END W2MID[3]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2114 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.512 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 7.80646 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 38.1791 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 13.620000 40.020000 14.000000 ;
    END
  END W2MID[2]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 5.93811 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 13.7145 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 12.400000 40.020000 12.780000 ;
    END
  END W2MID[1]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 39.320000 10.570000 40.020000 10.950000 ;
    END
  END W2MID[0]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 39.320000 33.140000 40.020000 33.520000 ;
    END
  END W2END[7]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.92 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 5.22364 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 23.6256 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 31.310000 40.020000 31.690000 ;
    END
  END W2END[6]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 3.74882 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 17.5448 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 30.090000 40.020000 30.470000 ;
    END
  END W2END[5]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 39.320000 28.870000 40.020000 29.250000 ;
    END
  END W2END[4]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 39.320000 27.040000 40.020000 27.420000 ;
    END
  END W2END[3]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3726 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.8398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 31.616 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 10.1537 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 53.2754 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 25.820000 40.020000 26.200000 ;
    END
  END W2END[2]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9544 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.752 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 7.07811 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 35.2444 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 23.990000 40.020000 24.370000 ;
    END
  END W2END[1]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 39.320000 22.770000 40.020000 23.150000 ;
    END
  END W2END[0]
  PIN WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9654 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.144 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 13.9398 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 70.0067 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 56.930000 40.020000 57.310000 ;
    END
  END WW4END[15]
  PIN WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 8.23286 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 40.0889 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 55.100000 40.020000 55.480000 ;
    END
  END WW4END[14]
  PIN WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 10.3589 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 50.3125 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 53.880000 40.020000 54.260000 ;
    END
  END WW4END[13]
  PIN WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2006 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.3668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 55.76 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 20.1981 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 105.837 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 52.660000 40.020000 53.040000 ;
    END
  END WW4END[12]
  PIN WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 7.51098 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 35.93 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 50.830000 40.020000 51.210000 ;
    END
  END WW4END[11]
  PIN WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0224 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 8.14343 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 39.7037 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 49.610000 40.020000 49.990000 ;
    END
  END WW4END[10]
  PIN WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 2.61212 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 11.6875 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 47.780000 40.020000 48.160000 ;
    END
  END WW4END[9]
  PIN WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.896 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 6.60458 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 32.2155 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 46.560000 40.020000 46.940000 ;
    END
  END WW4END[8]
  PIN WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 5.84875 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 27.7616 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 44.730000 40.020000 45.110000 ;
    END
  END WW4END[7]
  PIN WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.536 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 12.8427 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 64.9751 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 43.510000 40.020000 43.890000 ;
    END
  END WW4END[6]
  PIN WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 5.96997 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 28.6505 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 42.290000 40.020000 42.670000 ;
    END
  END WW4END[5]
  PIN WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8694 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.632 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 2.52848 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 11.7266 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 40.460000 40.020000 40.840000 ;
    END
  END WW4END[4]
  PIN WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 7.27475 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 36.0418 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 39.240000 40.020000 39.620000 ;
    END
  END WW4END[3]
  PIN WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 4.63906 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 21.8222 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 37.410000 40.020000 37.790000 ;
    END
  END WW4END[2]
  PIN WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 5.35232 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 25.2956 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 36.190000 40.020000 36.570000 ;
    END
  END WW4END[1]
  PIN WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 2.25939 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 9.87205 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 34.360000 40.020000 34.740000 ;
    END
  END WW4END[0]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.488 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 28.4329 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 134.575 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.477381 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 74.620000 40.020000 75.000000 ;
    END
  END W6END[11]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 41.8655 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 198.105 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 73.400000 40.020000 73.780000 ;
    END
  END W6END[10]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5964 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.176 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 31.1274 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 148.714 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.477381 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 71.570000 40.020000 71.950000 ;
    END
  END W6END[9]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.44 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 40.856 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 197.613 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 70.350000 40.020000 70.730000 ;
    END
  END W6END[8]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4834 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 36.9044 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 180.095 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.477381 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 68.520000 40.020000 68.900000 ;
    END
  END W6END[7]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 21.8357 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 96.7163 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 67.300000 40.020000 67.680000 ;
    END
  END W6END[6]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.104 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 52.2373 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 257.097 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 66.080000 40.020000 66.460000 ;
    END
  END W6END[5]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.696 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 53.9619 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 264.915 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 64.250000 40.020000 64.630000 ;
    END
  END W6END[4]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0074 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.368 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 49.2734 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 240.427 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 63.030000 40.020000 63.410000 ;
    END
  END W6END[3]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 41.0909 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 194.915 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 61.200000 40.020000 61.580000 ;
    END
  END W6END[2]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 19.4409 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 85.496 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.477381 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 59.980000 40.020000 60.360000 ;
    END
  END W6END[1]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.192 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 52.256 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 257.28 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 58.150000 40.020000 58.530000 ;
    END
  END W6END[0]
  PIN OPA_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6184 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.96 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 49.077 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 239.772 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 64.250000 0.700000 64.630000 ;
    END
  END OPA_I0
  PIN OPA_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5486 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.8178 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 52.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 47.9365 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 246.698 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 67.910000 0.700000 68.290000 ;
    END
  END OPA_I1
  PIN OPA_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8614 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.256 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 33.2798 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 159.839 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.566667 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 71.570000 0.700000 71.950000 ;
    END
  END OPA_I2
  PIN OPA_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6074 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.568 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 47.1766 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 230.736 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 75.230000 0.700000 75.610000 ;
    END
  END OPA_I3
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8029 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.608 LAYER met3  ;
    ANTENNAMAXAREACAR 2.33459 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 11.0039 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.0386502 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 0.000000 5.480000 0.700000 ;
    END
  END UserCLK
  PIN OPB_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 44.6595 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 210.272 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 49.000000 0.700000 49.380000 ;
    END
  END OPB_I0
  PIN OPB_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.5368 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 62.3536 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 315.819 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 53.270000 0.700000 53.650000 ;
    END
  END OPB_I1
  PIN OPB_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5434 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.56 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 45.1056 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 220.796 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.566667 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 56.930000 0.700000 57.310000 ;
    END
  END OPB_I2
  PIN OPB_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 25.6163 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 117.597 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 60.590000 0.700000 60.970000 ;
    END
  END OPB_I3
  PIN RES0_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 34.360000 0.700000 34.740000 ;
    END
  END RES0_O0
  PIN RES0_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 38.020000 0.700000 38.400000 ;
    END
  END RES0_O1
  PIN RES0_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 41.680000 0.700000 42.060000 ;
    END
  END RES0_O2
  PIN RES0_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 45.340000 0.700000 45.720000 ;
    END
  END RES0_O3
  PIN RES1_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 19.720000 0.700000 20.100000 ;
    END
  END RES1_O0
  PIN RES1_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 23.380000 0.700000 23.760000 ;
    END
  END RES1_O1
  PIN RES1_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 27.040000 0.700000 27.420000 ;
    END
  END RES1_O2
  PIN RES1_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 30.700000 0.700000 31.080000 ;
    END
  END RES1_O3
  PIN RES2_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 5.080000 0.700000 5.460000 ;
    END
  END RES2_O0
  PIN RES2_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.2644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.072 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 8.740000 0.700000 9.120000 ;
    END
  END RES2_O1
  PIN RES2_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2476 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.3448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 92.976 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 12.400000 0.700000 12.780000 ;
    END
  END RES2_O2
  PIN RES2_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 16.060000 0.700000 16.440000 ;
    END
  END RES2_O3
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 4.5209 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.8898 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.216 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 199.560000 5.480000 200.260000 ;
    END
  END UserCLKo
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.3224 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 32.9344 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 163.618 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 193.570000 0.700000 193.950000 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 6.07275 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 27.1817 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.25109 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 189.910000 0.700000 190.290000 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 12.6227 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 59.566 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 186.250000 0.700000 186.630000 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.96 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 19.8166 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 96.556 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 182.590000 0.700000 182.970000 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 4.39611 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 20.4885 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 178.930000 0.700000 179.310000 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6935 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.352 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 7.57246 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 36.8916 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.0488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 54.064 LAYER met4  ;
    ANTENNAGATEAREA 0.9015 LAYER met4  ;
    ANTENNAMAXAREACAR 19.7046 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 103.021 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 175.270000 0.700000 175.650000 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3213 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.704 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 15.2786 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 74.3897 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 171.610000 0.700000 171.990000 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 5.8367 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 25.8328 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.25109 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 167.950000 0.700000 168.330000 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.176 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 15.2871 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 78.9239 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 23.9088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 127.984 LAYER met4  ;
    ANTENNAGATEAREA 0.9015 LAYER met4  ;
    ANTENNAMAXAREACAR 50.6815 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 266.462 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 164.290000 0.700000 164.670000 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7056 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.088 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.9167 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 106.688 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met4  ;
    ANTENNAMAXAREACAR 59.8985 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 311.543 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 160.630000 0.700000 161.010000 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.816 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 18.6317 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 92.4276 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 156.970000 0.700000 157.350000 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 19.8108 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 95.5174 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 153.310000 0.700000 153.690000 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4493 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.72 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 24.6398 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 119.491 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 149.650000 0.700000 150.030000 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.96 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 16.6475 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 80.7216 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 145.380000 0.700000 145.760000 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0224 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 36.722 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 179.823 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.50915 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 141.720000 0.700000 142.100000 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1634 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 17.7356 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 86.4559 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 138.060000 0.700000 138.440000 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8283 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.408 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 21.9637 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 107.811 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 134.400000 0.700000 134.780000 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.432 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 14.2039 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 68.5072 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 130.740000 0.700000 131.120000 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.216 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 59.3138 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 306.204 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.4388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.144 LAYER met4  ;
    ANTENNAGATEAREA 0.9015 LAYER met4  ;
    ANTENNAMAXAREACAR 67.5654 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 350.735 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 127.080000 0.700000 127.460000 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3506 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.7907 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 58.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met4  ;
    ANTENNAMAXAREACAR 18.6653 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 96.7921 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 123.420000 0.700000 123.800000 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.1578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 16.6003 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 87.5071 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 119.760000 0.700000 120.140000 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 8.71232 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 42.0956 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 116.100000 0.700000 116.480000 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.68 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 13.772 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 70.1387 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 112.440000 0.700000 112.820000 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 11.2265 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 56.563 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 108.780000 0.700000 109.160000 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 5.76465 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 26.2047 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 105.120000 0.700000 105.500000 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6836 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.8048 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 42.096 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 14.4998 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 76.6182 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 101.460000 0.700000 101.840000 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.1578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 14.3906 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 75.868 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 97.190000 0.700000 97.570000 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 6.2767 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 29.3145 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 93.530000 0.700000 93.910000 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5754 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.064 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 5.77798 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 26.4256 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 89.870000 0.700000 90.250000 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7428 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.432 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 11.2703 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 58.637 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 86.210000 0.700000 86.590000 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7536 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.1378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 91.872 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 24.3801 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 129.592 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 82.550000 0.700000 82.930000 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5774 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.408 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 13.6178 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 67.3805 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 78.890000 0.700000 79.270000 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 194.180000 40.020000 194.560000 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 192.350000 40.020000 192.730000 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 191.130000 40.020000 191.510000 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.4474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.048 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 189.300000 40.020000 189.680000 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.1034 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.88 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 188.080000 40.020000 188.460000 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.9884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 186.250000 40.020000 186.630000 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 185.030000 40.020000 185.410000 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 183.200000 40.020000 183.580000 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 181.980000 40.020000 182.360000 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 180.760000 40.020000 181.140000 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 178.930000 40.020000 179.310000 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.2644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.072 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 177.710000 40.020000 178.090000 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 175.880000 40.020000 176.260000 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.7824 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.168 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 174.660000 40.020000 175.040000 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 172.830000 40.020000 173.210000 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 171.610000 40.020000 171.990000 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 169.780000 40.020000 170.160000 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 168.560000 40.020000 168.940000 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 167.340000 40.020000 167.720000 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 165.510000 40.020000 165.890000 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6146 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.6088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 30.384 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 164.290000 40.020000 164.670000 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9026 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.8158 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 31.488 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 162.460000 40.020000 162.840000 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 161.240000 40.020000 161.620000 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 159.410000 40.020000 159.790000 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7594 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.712 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 158.190000 40.020000 158.570000 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.712 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 156.360000 40.020000 156.740000 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 155.140000 40.020000 155.520000 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 153.920000 40.020000 154.300000 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.6214 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.976 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 152.090000 40.020000 152.470000 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.4724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.848 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 150.870000 40.020000 151.250000 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 149.040000 40.020000 149.420000 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3726 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.9748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.336 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 147.820000 40.020000 148.200000 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.8396 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 12.9125 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 34.540000 0.000000 34.920000 0.700000 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.5978 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 92.645 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 25.5749 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 126.176 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 32.700000 0.000000 33.080000 0.700000 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.4818 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 147.04 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 44.1733 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 233.09 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 31.320000 0.000000 31.700000 0.700000 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8277 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.9775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 39.3288 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 210.224 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 53.9467 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 287.442 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 29.940000 0.000000 30.320000 0.700000 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.529 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 97.419 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 28.2187 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 139.554 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 28.560000 0.000000 28.940000 0.700000 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7609 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 39.3288 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 210.224 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 54.2432 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 289.014 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 27.180000 0.000000 27.560000 0.700000 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8029 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.3658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 221.088 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 58.8136 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 312.924 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 25.340000 0.000000 25.720000 0.700000 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1087 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.3825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.0828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 176.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 48.4541 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 258.083 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 23.960000 0.000000 24.340000 0.700000 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.2562 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 96.173 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 26.4617 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 130.927 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 22.580000 0.000000 22.960000 0.700000 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2795 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.2365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 40.2438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 215.104 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 57.5692 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 306.726 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 21.200000 0.000000 21.580000 0.700000 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 46.2588 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 247.184 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 63.953 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 340.57 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 19.360000 0.000000 19.740000 0.700000 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.8853 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.1475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.299 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.1678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 172.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 48.2062 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 255.789 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 17.980000 0.000000 18.360000 0.700000 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 46.4658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 248.288 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 63.8333 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 340.269 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 16.600000 0.000000 16.980000 0.700000 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7175 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.1358 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.528 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 40.4669 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 208.048 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 15.220000 0.000000 15.600000 0.700000 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1766 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.775 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.53481 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.2431 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 13.840000 0.000000 14.220000 0.700000 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.7328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 73.712 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 45.1314 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 232.046 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 12.460000 0.000000 12.840000 0.700000 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 47.9058 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 255.968 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 65.503 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 349.051 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 10.620000 0.000000 11.000000 0.700000 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1445 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.1608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 241.328 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 62.0541 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 330.459 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 9.240000 0.000000 9.620000 0.700000 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.01872 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.8081 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 7.860000 0.000000 8.240000 0.700000 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.3116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 119.476 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3765 LAYER met2  ;
    ANTENNAMAXAREACAR 18.8229 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 88.5135 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.46478 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 6.480000 0.000000 6.860000 0.700000 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7482 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.633 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 34.540000 199.560000 34.920000 200.260000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4021 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.8438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.304 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 32.700000 199.560000 33.080000 200.260000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8897 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.3948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.576 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 31.320000 199.560000 31.700000 200.260000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.2578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 76.512 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 29.940000 199.560000 30.320000 200.260000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.8458 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.121 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 28.560000 199.560000 28.940000 200.260000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4913 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.2955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8088 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.784 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 27.180000 199.560000 27.560000 200.260000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.1598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.656 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 25.340000 199.560000 25.720000 200.260000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.2968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 108.72 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 23.960000 199.560000 24.340000 200.260000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.3974 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.879 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 22.580000 199.560000 22.960000 200.260000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.3034 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.409 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 21.200000 199.560000 21.580000 200.260000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.0014 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.899 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 19.360000 199.560000 19.740000 200.260000 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.4388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.144 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 17.980000 199.560000 18.360000 200.260000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.5246 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.515 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 16.600000 199.560000 16.980000 200.260000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.9562 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.673 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 15.220000 199.560000 15.600000 200.260000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.8614 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.199 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 13.840000 199.560000 14.220000 200.260000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.9638 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.593 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 12.460000 199.560000 12.840000 200.260000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.5618 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.701 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 10.620000 199.560000 11.000000 200.260000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.0514 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.149 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 9.240000 199.560000 9.620000 200.260000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.259 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.187 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 7.860000 199.560000 8.240000 200.260000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.4498 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.141 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 6.480000 199.560000 6.860000 200.260000 ;
    END
  END FrameStrobe_O[0]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 38.820000 195.020000 40.020000 196.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 195.020000 1.200000 196.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.820000 2.850000 40.020000 4.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 1.200000 4.050000 ;
    END
    PORT
      LAYER met4 ;
        RECT 35.990000 199.060000 37.190000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 35.990000 0.000000 37.190000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 199.060000 4.030000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 0.000000 4.030000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 40.020000 4.050000 ;
        RECT 0.000000 195.020000 40.020000 196.220000 ;
        RECT 2.830000 10.300000 4.030000 10.780000 ;
        RECT 2.830000 4.860000 4.030000 5.340000 ;
        RECT 7.060000 10.300000 8.260000 10.780000 ;
        RECT 7.060000 4.860000 8.260000 5.340000 ;
        RECT 7.060000 21.180000 8.260000 21.660000 ;
        RECT 7.060000 15.740000 8.260000 16.220000 ;
        RECT 2.830000 21.180000 4.030000 21.660000 ;
        RECT 2.830000 15.740000 4.030000 16.220000 ;
        RECT 2.830000 37.500000 4.030000 37.980000 ;
        RECT 7.060000 37.500000 8.260000 37.980000 ;
        RECT 2.830000 32.060000 4.030000 32.540000 ;
        RECT 2.830000 26.620000 4.030000 27.100000 ;
        RECT 7.060000 32.060000 8.260000 32.540000 ;
        RECT 7.060000 26.620000 8.260000 27.100000 ;
        RECT 2.830000 48.380000 4.030000 48.860000 ;
        RECT 2.830000 42.940000 4.030000 43.420000 ;
        RECT 7.060000 48.380000 8.260000 48.860000 ;
        RECT 7.060000 42.940000 8.260000 43.420000 ;
        RECT 7.060000 59.260000 8.260000 59.740000 ;
        RECT 7.060000 53.820000 8.260000 54.300000 ;
        RECT 2.830000 59.260000 4.030000 59.740000 ;
        RECT 2.830000 53.820000 4.030000 54.300000 ;
        RECT 2.830000 70.140000 4.030000 70.620000 ;
        RECT 2.830000 64.700000 4.030000 65.180000 ;
        RECT 7.060000 70.140000 8.260000 70.620000 ;
        RECT 7.060000 64.700000 8.260000 65.180000 ;
        RECT 7.060000 86.460000 8.260000 86.940000 ;
        RECT 7.060000 81.020000 8.260000 81.500000 ;
        RECT 7.060000 75.580000 8.260000 76.060000 ;
        RECT 2.830000 86.460000 4.030000 86.940000 ;
        RECT 2.830000 81.020000 4.030000 81.500000 ;
        RECT 2.830000 75.580000 4.030000 76.060000 ;
        RECT 2.830000 97.340000 4.030000 97.820000 ;
        RECT 2.830000 91.900000 4.030000 92.380000 ;
        RECT 7.060000 97.340000 8.260000 97.820000 ;
        RECT 7.060000 91.900000 8.260000 92.380000 ;
        RECT 35.990000 10.300000 37.190000 10.780000 ;
        RECT 35.990000 4.860000 37.190000 5.340000 ;
        RECT 35.990000 21.180000 37.190000 21.660000 ;
        RECT 35.990000 15.740000 37.190000 16.220000 ;
        RECT 35.990000 37.500000 37.190000 37.980000 ;
        RECT 35.990000 32.060000 37.190000 32.540000 ;
        RECT 35.990000 26.620000 37.190000 27.100000 ;
        RECT 35.990000 48.380000 37.190000 48.860000 ;
        RECT 35.990000 42.940000 37.190000 43.420000 ;
        RECT 35.990000 59.260000 37.190000 59.740000 ;
        RECT 35.990000 53.820000 37.190000 54.300000 ;
        RECT 35.990000 70.140000 37.190000 70.620000 ;
        RECT 35.990000 64.700000 37.190000 65.180000 ;
        RECT 35.990000 86.460000 37.190000 86.940000 ;
        RECT 35.990000 81.020000 37.190000 81.500000 ;
        RECT 35.990000 75.580000 37.190000 76.060000 ;
        RECT 35.990000 97.340000 37.190000 97.820000 ;
        RECT 35.990000 91.900000 37.190000 92.380000 ;
        RECT 2.830000 108.220000 4.030000 108.700000 ;
        RECT 2.830000 102.780000 4.030000 103.260000 ;
        RECT 7.060000 108.220000 8.260000 108.700000 ;
        RECT 7.060000 102.780000 8.260000 103.260000 ;
        RECT 7.060000 124.540000 8.260000 125.020000 ;
        RECT 7.060000 119.100000 8.260000 119.580000 ;
        RECT 7.060000 113.660000 8.260000 114.140000 ;
        RECT 2.830000 124.540000 4.030000 125.020000 ;
        RECT 2.830000 119.100000 4.030000 119.580000 ;
        RECT 2.830000 113.660000 4.030000 114.140000 ;
        RECT 2.830000 135.420000 4.030000 135.900000 ;
        RECT 2.830000 129.980000 4.030000 130.460000 ;
        RECT 7.060000 135.420000 8.260000 135.900000 ;
        RECT 7.060000 129.980000 8.260000 130.460000 ;
        RECT 7.060000 146.300000 8.260000 146.780000 ;
        RECT 7.060000 140.860000 8.260000 141.340000 ;
        RECT 2.830000 146.300000 4.030000 146.780000 ;
        RECT 2.830000 140.860000 4.030000 141.340000 ;
        RECT 2.830000 162.620000 4.030000 163.100000 ;
        RECT 7.060000 162.620000 8.260000 163.100000 ;
        RECT 2.830000 157.180000 4.030000 157.660000 ;
        RECT 2.830000 151.740000 4.030000 152.220000 ;
        RECT 7.060000 157.180000 8.260000 157.660000 ;
        RECT 7.060000 151.740000 8.260000 152.220000 ;
        RECT 2.830000 173.500000 4.030000 173.980000 ;
        RECT 2.830000 168.060000 4.030000 168.540000 ;
        RECT 7.060000 173.500000 8.260000 173.980000 ;
        RECT 7.060000 168.060000 8.260000 168.540000 ;
        RECT 7.060000 184.380000 8.260000 184.860000 ;
        RECT 7.060000 178.940000 8.260000 179.420000 ;
        RECT 2.830000 184.380000 4.030000 184.860000 ;
        RECT 2.830000 178.940000 4.030000 179.420000 ;
        RECT 2.830000 189.820000 4.030000 190.300000 ;
        RECT 7.060000 189.820000 8.260000 190.300000 ;
        RECT 35.990000 108.220000 37.190000 108.700000 ;
        RECT 35.990000 102.780000 37.190000 103.260000 ;
        RECT 35.990000 124.540000 37.190000 125.020000 ;
        RECT 35.990000 119.100000 37.190000 119.580000 ;
        RECT 35.990000 113.660000 37.190000 114.140000 ;
        RECT 35.990000 135.420000 37.190000 135.900000 ;
        RECT 35.990000 129.980000 37.190000 130.460000 ;
        RECT 35.990000 146.300000 37.190000 146.780000 ;
        RECT 35.990000 140.860000 37.190000 141.340000 ;
        RECT 35.990000 162.620000 37.190000 163.100000 ;
        RECT 35.990000 157.180000 37.190000 157.660000 ;
        RECT 35.990000 151.740000 37.190000 152.220000 ;
        RECT 35.990000 173.500000 37.190000 173.980000 ;
        RECT 35.990000 168.060000 37.190000 168.540000 ;
        RECT 35.990000 178.940000 37.190000 179.420000 ;
        RECT 35.990000 184.380000 37.190000 184.860000 ;
        RECT 35.990000 189.820000 37.190000 190.300000 ;
      LAYER met4 ;
        RECT 7.060000 2.850000 8.260000 196.220000 ;
        RECT 35.990000 0.000000 37.190000 200.260000 ;
        RECT 2.830000 0.000000 4.030000 200.260000 ;
    END
# end of P/G power stripe data as pin

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 38.820000 196.820000 40.020000 198.020000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 196.820000 1.200000 198.020000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.820000 1.050000 40.020000 2.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 1.200000 2.250000 ;
    END
    PORT
      LAYER met4 ;
        RECT 37.790000 199.060000 38.990000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 37.790000 0.000000 38.990000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 199.060000 2.230000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 0.000000 2.230000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 40.020000 2.250000 ;
        RECT 0.000000 196.820000 40.020000 198.020000 ;
        RECT 37.790000 100.060000 38.990000 100.540000 ;
        RECT 1.030000 100.060000 2.230000 100.540000 ;
        RECT 4.895000 100.060000 6.260000 100.540000 ;
        RECT 1.030000 7.580000 2.230000 8.060000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
        RECT 1.030000 13.020000 2.230000 13.500000 ;
        RECT 1.030000 18.460000 2.230000 18.940000 ;
        RECT 1.030000 23.900000 2.230000 24.380000 ;
        RECT 1.030000 34.780000 2.230000 35.260000 ;
        RECT 1.030000 29.340000 2.230000 29.820000 ;
        RECT 4.895000 34.780000 6.260000 35.260000 ;
        RECT 4.895000 29.340000 6.260000 29.820000 ;
        RECT 1.030000 45.660000 2.230000 46.140000 ;
        RECT 1.030000 40.220000 2.230000 40.700000 ;
        RECT 4.895000 45.660000 6.260000 46.140000 ;
        RECT 4.895000 40.220000 6.260000 40.700000 ;
        RECT 1.030000 51.100000 2.230000 51.580000 ;
        RECT 4.895000 51.100000 6.260000 51.580000 ;
        RECT 4.895000 56.540000 6.260000 57.020000 ;
        RECT 4.895000 61.980000 6.260000 62.460000 ;
        RECT 1.030000 56.540000 2.230000 57.020000 ;
        RECT 1.030000 61.980000 2.230000 62.460000 ;
        RECT 1.030000 72.860000 2.230000 73.340000 ;
        RECT 1.030000 67.420000 2.230000 67.900000 ;
        RECT 4.895000 72.860000 6.260000 73.340000 ;
        RECT 4.895000 67.420000 6.260000 67.900000 ;
        RECT 4.895000 78.300000 6.260000 78.780000 ;
        RECT 4.895000 83.740000 6.260000 84.220000 ;
        RECT 1.030000 78.300000 2.230000 78.780000 ;
        RECT 1.030000 83.740000 2.230000 84.220000 ;
        RECT 1.030000 94.620000 2.230000 95.100000 ;
        RECT 1.030000 89.180000 2.230000 89.660000 ;
        RECT 4.895000 94.620000 6.260000 95.100000 ;
        RECT 4.895000 89.180000 6.260000 89.660000 ;
        RECT 37.790000 7.580000 38.990000 8.060000 ;
        RECT 37.790000 23.900000 38.990000 24.380000 ;
        RECT 37.790000 18.460000 38.990000 18.940000 ;
        RECT 37.790000 13.020000 38.990000 13.500000 ;
        RECT 37.790000 29.340000 38.990000 29.820000 ;
        RECT 37.790000 34.780000 38.990000 35.260000 ;
        RECT 37.790000 45.660000 38.990000 46.140000 ;
        RECT 37.790000 40.220000 38.990000 40.700000 ;
        RECT 37.790000 61.980000 38.990000 62.460000 ;
        RECT 37.790000 56.540000 38.990000 57.020000 ;
        RECT 37.790000 51.100000 38.990000 51.580000 ;
        RECT 37.790000 72.860000 38.990000 73.340000 ;
        RECT 37.790000 67.420000 38.990000 67.900000 ;
        RECT 37.790000 83.740000 38.990000 84.220000 ;
        RECT 37.790000 78.300000 38.990000 78.780000 ;
        RECT 37.790000 94.620000 38.990000 95.100000 ;
        RECT 37.790000 89.180000 38.990000 89.660000 ;
        RECT 1.030000 110.940000 2.230000 111.420000 ;
        RECT 1.030000 105.500000 2.230000 105.980000 ;
        RECT 4.895000 110.940000 6.260000 111.420000 ;
        RECT 4.895000 105.500000 6.260000 105.980000 ;
        RECT 4.895000 121.820000 6.260000 122.300000 ;
        RECT 4.895000 116.380000 6.260000 116.860000 ;
        RECT 1.030000 116.380000 2.230000 116.860000 ;
        RECT 1.030000 121.820000 2.230000 122.300000 ;
        RECT 1.030000 132.700000 2.230000 133.180000 ;
        RECT 4.895000 132.700000 6.260000 133.180000 ;
        RECT 4.895000 127.260000 6.260000 127.740000 ;
        RECT 1.030000 127.260000 2.230000 127.740000 ;
        RECT 4.895000 138.140000 6.260000 138.620000 ;
        RECT 4.895000 143.580000 6.260000 144.060000 ;
        RECT 4.895000 149.020000 6.260000 149.500000 ;
        RECT 1.030000 138.140000 2.230000 138.620000 ;
        RECT 1.030000 143.580000 2.230000 144.060000 ;
        RECT 1.030000 149.020000 2.230000 149.500000 ;
        RECT 1.030000 159.900000 2.230000 160.380000 ;
        RECT 1.030000 154.460000 2.230000 154.940000 ;
        RECT 4.895000 159.900000 6.260000 160.380000 ;
        RECT 4.895000 154.460000 6.260000 154.940000 ;
        RECT 1.030000 170.780000 2.230000 171.260000 ;
        RECT 1.030000 165.340000 2.230000 165.820000 ;
        RECT 4.895000 170.780000 6.260000 171.260000 ;
        RECT 4.895000 165.340000 6.260000 165.820000 ;
        RECT 4.895000 176.220000 6.260000 176.700000 ;
        RECT 4.895000 181.660000 6.260000 182.140000 ;
        RECT 4.895000 187.100000 6.260000 187.580000 ;
        RECT 1.030000 176.220000 2.230000 176.700000 ;
        RECT 1.030000 181.660000 2.230000 182.140000 ;
        RECT 1.030000 187.100000 2.230000 187.580000 ;
        RECT 1.030000 192.540000 2.230000 193.020000 ;
        RECT 4.895000 192.540000 6.260000 193.020000 ;
        RECT 37.790000 110.940000 38.990000 111.420000 ;
        RECT 37.790000 105.500000 38.990000 105.980000 ;
        RECT 37.790000 116.380000 38.990000 116.860000 ;
        RECT 37.790000 121.820000 38.990000 122.300000 ;
        RECT 37.790000 132.700000 38.990000 133.180000 ;
        RECT 37.790000 127.260000 38.990000 127.740000 ;
        RECT 37.790000 149.020000 38.990000 149.500000 ;
        RECT 37.790000 143.580000 38.990000 144.060000 ;
        RECT 37.790000 138.140000 38.990000 138.620000 ;
        RECT 37.790000 159.900000 38.990000 160.380000 ;
        RECT 37.790000 154.460000 38.990000 154.940000 ;
        RECT 37.790000 170.780000 38.990000 171.260000 ;
        RECT 37.790000 165.340000 38.990000 165.820000 ;
        RECT 37.790000 181.660000 38.990000 182.140000 ;
        RECT 37.790000 176.220000 38.990000 176.700000 ;
        RECT 37.790000 187.100000 38.990000 187.580000 ;
        RECT 37.790000 192.540000 38.990000 193.020000 ;
      LAYER met4 ;
        RECT 5.060000 1.050000 6.260000 198.020000 ;
        RECT 37.790000 0.000000 38.990000 200.260000 ;
        RECT 1.030000 0.000000 2.230000 200.260000 ;
        RECT 4.895000 100.060000 6.260000 100.540000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
        RECT 4.895000 34.780000 6.260000 35.260000 ;
        RECT 4.895000 29.340000 6.260000 29.820000 ;
        RECT 4.895000 45.660000 6.260000 46.140000 ;
        RECT 4.895000 40.220000 6.260000 40.700000 ;
        RECT 4.895000 51.100000 6.260000 51.580000 ;
        RECT 4.895000 56.540000 6.260000 57.020000 ;
        RECT 4.895000 61.980000 6.260000 62.460000 ;
        RECT 4.895000 72.860000 6.260000 73.340000 ;
        RECT 4.895000 67.420000 6.260000 67.900000 ;
        RECT 4.895000 78.300000 6.260000 78.780000 ;
        RECT 4.895000 83.740000 6.260000 84.220000 ;
        RECT 4.895000 94.620000 6.260000 95.100000 ;
        RECT 4.895000 89.180000 6.260000 89.660000 ;
        RECT 4.895000 110.940000 6.260000 111.420000 ;
        RECT 4.895000 105.500000 6.260000 105.980000 ;
        RECT 4.895000 121.820000 6.260000 122.300000 ;
        RECT 4.895000 116.380000 6.260000 116.860000 ;
        RECT 4.895000 132.700000 6.260000 133.180000 ;
        RECT 4.895000 127.260000 6.260000 127.740000 ;
        RECT 4.895000 138.140000 6.260000 138.620000 ;
        RECT 4.895000 143.580000 6.260000 144.060000 ;
        RECT 4.895000 149.020000 6.260000 149.500000 ;
        RECT 4.895000 159.900000 6.260000 160.380000 ;
        RECT 4.895000 154.460000 6.260000 154.940000 ;
        RECT 4.895000 170.780000 6.260000 171.260000 ;
        RECT 4.895000 165.340000 6.260000 165.820000 ;
        RECT 4.895000 176.220000 6.260000 176.700000 ;
        RECT 4.895000 181.660000 6.260000 182.140000 ;
        RECT 4.895000 187.100000 6.260000 187.580000 ;
        RECT 4.895000 192.540000 6.260000 193.020000 ;
    END
# end of P/G power stripe data as pin

  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 40.020000 200.260000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 40.020000 200.260000 ;
    LAYER met2 ;
      RECT 35.060000 199.420000 40.020000 200.260000 ;
      RECT 33.220000 199.420000 34.400000 200.260000 ;
      RECT 31.840000 199.420000 32.560000 200.260000 ;
      RECT 30.460000 199.420000 31.180000 200.260000 ;
      RECT 29.080000 199.420000 29.800000 200.260000 ;
      RECT 27.700000 199.420000 28.420000 200.260000 ;
      RECT 25.860000 199.420000 27.040000 200.260000 ;
      RECT 24.480000 199.420000 25.200000 200.260000 ;
      RECT 23.100000 199.420000 23.820000 200.260000 ;
      RECT 21.720000 199.420000 22.440000 200.260000 ;
      RECT 19.880000 199.420000 21.060000 200.260000 ;
      RECT 18.500000 199.420000 19.220000 200.260000 ;
      RECT 17.120000 199.420000 17.840000 200.260000 ;
      RECT 15.740000 199.420000 16.460000 200.260000 ;
      RECT 14.360000 199.420000 15.080000 200.260000 ;
      RECT 12.980000 199.420000 13.700000 200.260000 ;
      RECT 11.140000 199.420000 12.320000 200.260000 ;
      RECT 9.760000 199.420000 10.480000 200.260000 ;
      RECT 8.380000 199.420000 9.100000 200.260000 ;
      RECT 7.000000 199.420000 7.720000 200.260000 ;
      RECT 5.620000 199.420000 6.340000 200.260000 ;
      RECT 0.000000 199.420000 4.960000 200.260000 ;
      RECT 0.000000 0.840000 40.020000 199.420000 ;
      RECT 35.060000 0.000000 40.020000 0.840000 ;
      RECT 33.220000 0.000000 34.400000 0.840000 ;
      RECT 31.840000 0.000000 32.560000 0.840000 ;
      RECT 30.460000 0.000000 31.180000 0.840000 ;
      RECT 29.080000 0.000000 29.800000 0.840000 ;
      RECT 27.700000 0.000000 28.420000 0.840000 ;
      RECT 25.860000 0.000000 27.040000 0.840000 ;
      RECT 24.480000 0.000000 25.200000 0.840000 ;
      RECT 23.100000 0.000000 23.820000 0.840000 ;
      RECT 21.720000 0.000000 22.440000 0.840000 ;
      RECT 19.880000 0.000000 21.060000 0.840000 ;
      RECT 18.500000 0.000000 19.220000 0.840000 ;
      RECT 17.120000 0.000000 17.840000 0.840000 ;
      RECT 15.740000 0.000000 16.460000 0.840000 ;
      RECT 14.360000 0.000000 15.080000 0.840000 ;
      RECT 12.980000 0.000000 13.700000 0.840000 ;
      RECT 11.140000 0.000000 12.320000 0.840000 ;
      RECT 9.760000 0.000000 10.480000 0.840000 ;
      RECT 8.380000 0.000000 9.100000 0.840000 ;
      RECT 7.000000 0.000000 7.720000 0.840000 ;
      RECT 5.620000 0.000000 6.340000 0.840000 ;
      RECT 0.000000 0.000000 4.960000 0.840000 ;
    LAYER met3 ;
      RECT 0.000000 198.320000 40.020000 200.260000 ;
      RECT 0.000000 194.250000 39.020000 194.720000 ;
      RECT 1.000000 193.880000 39.020000 194.250000 ;
      RECT 1.000000 193.320000 40.020000 193.880000 ;
      RECT 39.290000 193.030000 40.020000 193.320000 ;
      RECT 6.560000 192.240000 37.490000 193.320000 ;
      RECT 2.530000 192.240000 4.595000 193.320000 ;
      RECT 0.000000 192.240000 0.730000 193.270000 ;
      RECT 0.000000 192.050000 39.020000 192.240000 ;
      RECT 0.000000 191.810000 40.020000 192.050000 ;
      RECT 0.000000 190.830000 39.020000 191.810000 ;
      RECT 0.000000 190.600000 40.020000 190.830000 ;
      RECT 0.000000 190.590000 2.530000 190.600000 ;
      RECT 37.490000 189.980000 40.020000 190.600000 ;
      RECT 1.000000 189.610000 2.530000 190.590000 ;
      RECT 37.490000 189.520000 39.020000 189.980000 ;
      RECT 8.560000 189.520000 35.690000 190.600000 ;
      RECT 4.330000 189.520000 6.760000 190.600000 ;
      RECT 0.000000 189.520000 2.530000 189.610000 ;
      RECT 0.000000 189.000000 39.020000 189.520000 ;
      RECT 0.000000 188.760000 40.020000 189.000000 ;
      RECT 0.000000 187.880000 39.020000 188.760000 ;
      RECT 39.290000 186.930000 40.020000 187.780000 ;
      RECT 0.000000 186.930000 0.730000 187.880000 ;
      RECT 6.560000 186.800000 37.490000 187.880000 ;
      RECT 2.530000 186.800000 4.595000 187.880000 ;
      RECT 1.000000 185.950000 39.020000 186.800000 ;
      RECT 0.000000 185.710000 40.020000 185.950000 ;
      RECT 0.000000 185.160000 39.020000 185.710000 ;
      RECT 37.490000 184.730000 39.020000 185.160000 ;
      RECT 37.490000 184.080000 40.020000 184.730000 ;
      RECT 8.560000 184.080000 35.690000 185.160000 ;
      RECT 4.330000 184.080000 6.760000 185.160000 ;
      RECT 0.000000 184.080000 2.530000 185.160000 ;
      RECT 0.000000 183.880000 40.020000 184.080000 ;
      RECT 0.000000 183.270000 39.020000 183.880000 ;
      RECT 1.000000 182.900000 39.020000 183.270000 ;
      RECT 1.000000 182.660000 40.020000 182.900000 ;
      RECT 1.000000 182.440000 39.020000 182.660000 ;
      RECT 39.290000 181.440000 40.020000 181.680000 ;
      RECT 6.560000 181.360000 37.490000 182.440000 ;
      RECT 2.530000 181.360000 4.595000 182.440000 ;
      RECT 0.000000 181.360000 0.730000 182.290000 ;
      RECT 0.000000 180.460000 39.020000 181.360000 ;
      RECT 0.000000 179.720000 40.020000 180.460000 ;
      RECT 37.490000 179.610000 40.020000 179.720000 ;
      RECT 0.000000 179.610000 2.530000 179.720000 ;
      RECT 37.490000 178.640000 39.020000 179.610000 ;
      RECT 8.560000 178.640000 35.690000 179.720000 ;
      RECT 4.330000 178.640000 6.760000 179.720000 ;
      RECT 1.000000 178.640000 2.530000 179.610000 ;
      RECT 1.000000 178.630000 39.020000 178.640000 ;
      RECT 0.000000 178.390000 40.020000 178.630000 ;
      RECT 0.000000 177.410000 39.020000 178.390000 ;
      RECT 0.000000 177.000000 40.020000 177.410000 ;
      RECT 39.290000 176.560000 40.020000 177.000000 ;
      RECT 0.000000 175.950000 0.730000 177.000000 ;
      RECT 6.560000 175.920000 37.490000 177.000000 ;
      RECT 2.530000 175.920000 4.595000 177.000000 ;
      RECT 1.000000 175.580000 39.020000 175.920000 ;
      RECT 1.000000 175.340000 40.020000 175.580000 ;
      RECT 1.000000 174.970000 39.020000 175.340000 ;
      RECT 0.000000 174.360000 39.020000 174.970000 ;
      RECT 0.000000 174.280000 40.020000 174.360000 ;
      RECT 37.490000 173.510000 40.020000 174.280000 ;
      RECT 37.490000 173.200000 39.020000 173.510000 ;
      RECT 8.560000 173.200000 35.690000 174.280000 ;
      RECT 4.330000 173.200000 6.760000 174.280000 ;
      RECT 0.000000 173.200000 2.530000 174.280000 ;
      RECT 0.000000 172.530000 39.020000 173.200000 ;
      RECT 0.000000 172.290000 40.020000 172.530000 ;
      RECT 1.000000 171.560000 39.020000 172.290000 ;
      RECT 39.290000 170.480000 40.020000 171.310000 ;
      RECT 6.560000 170.480000 37.490000 171.560000 ;
      RECT 2.530000 170.480000 4.595000 171.560000 ;
      RECT 0.000000 170.480000 0.730000 171.310000 ;
      RECT 0.000000 170.460000 40.020000 170.480000 ;
      RECT 0.000000 169.480000 39.020000 170.460000 ;
      RECT 0.000000 169.240000 40.020000 169.480000 ;
      RECT 0.000000 168.840000 39.020000 169.240000 ;
      RECT 0.000000 168.630000 2.530000 168.840000 ;
      RECT 37.490000 168.260000 39.020000 168.840000 ;
      RECT 37.490000 168.020000 40.020000 168.260000 ;
      RECT 37.490000 167.760000 39.020000 168.020000 ;
      RECT 8.560000 167.760000 35.690000 168.840000 ;
      RECT 4.330000 167.760000 6.760000 168.840000 ;
      RECT 1.000000 167.760000 2.530000 168.630000 ;
      RECT 1.000000 167.650000 39.020000 167.760000 ;
      RECT 0.000000 167.040000 39.020000 167.650000 ;
      RECT 0.000000 166.190000 40.020000 167.040000 ;
      RECT 0.000000 166.120000 39.020000 166.190000 ;
      RECT 39.290000 165.040000 40.020000 165.210000 ;
      RECT 6.560000 165.040000 37.490000 166.120000 ;
      RECT 2.530000 165.040000 4.595000 166.120000 ;
      RECT 0.000000 165.040000 0.730000 166.120000 ;
      RECT 0.000000 164.970000 40.020000 165.040000 ;
      RECT 1.000000 163.990000 39.020000 164.970000 ;
      RECT 0.000000 163.400000 40.020000 163.990000 ;
      RECT 37.490000 163.140000 40.020000 163.400000 ;
      RECT 37.490000 162.320000 39.020000 163.140000 ;
      RECT 8.560000 162.320000 35.690000 163.400000 ;
      RECT 4.330000 162.320000 6.760000 163.400000 ;
      RECT 0.000000 162.320000 2.530000 163.400000 ;
      RECT 0.000000 162.160000 39.020000 162.320000 ;
      RECT 0.000000 161.920000 40.020000 162.160000 ;
      RECT 0.000000 161.310000 39.020000 161.920000 ;
      RECT 1.000000 160.940000 39.020000 161.310000 ;
      RECT 1.000000 160.680000 40.020000 160.940000 ;
      RECT 39.290000 160.090000 40.020000 160.680000 ;
      RECT 6.560000 159.600000 37.490000 160.680000 ;
      RECT 2.530000 159.600000 4.595000 160.680000 ;
      RECT 0.000000 159.600000 0.730000 160.330000 ;
      RECT 0.000000 159.110000 39.020000 159.600000 ;
      RECT 0.000000 158.870000 40.020000 159.110000 ;
      RECT 0.000000 157.960000 39.020000 158.870000 ;
      RECT 37.490000 157.890000 39.020000 157.960000 ;
      RECT 0.000000 157.650000 2.530000 157.960000 ;
      RECT 37.490000 157.040000 40.020000 157.890000 ;
      RECT 37.490000 156.880000 39.020000 157.040000 ;
      RECT 8.560000 156.880000 35.690000 157.960000 ;
      RECT 4.330000 156.880000 6.760000 157.960000 ;
      RECT 1.000000 156.880000 2.530000 157.650000 ;
      RECT 1.000000 156.670000 39.020000 156.880000 ;
      RECT 0.000000 156.060000 39.020000 156.670000 ;
      RECT 0.000000 155.820000 40.020000 156.060000 ;
      RECT 0.000000 155.240000 39.020000 155.820000 ;
      RECT 39.290000 154.600000 40.020000 154.840000 ;
      RECT 6.560000 154.160000 37.490000 155.240000 ;
      RECT 2.530000 154.160000 4.595000 155.240000 ;
      RECT 0.000000 154.160000 0.730000 155.240000 ;
      RECT 0.000000 153.990000 39.020000 154.160000 ;
      RECT 1.000000 153.620000 39.020000 153.990000 ;
      RECT 1.000000 153.010000 40.020000 153.620000 ;
      RECT 0.000000 152.770000 40.020000 153.010000 ;
      RECT 0.000000 152.520000 39.020000 152.770000 ;
      RECT 37.490000 151.790000 39.020000 152.520000 ;
      RECT 37.490000 151.550000 40.020000 151.790000 ;
      RECT 37.490000 151.440000 39.020000 151.550000 ;
      RECT 8.560000 151.440000 35.690000 152.520000 ;
      RECT 4.330000 151.440000 6.760000 152.520000 ;
      RECT 0.000000 151.440000 2.530000 152.520000 ;
      RECT 0.000000 150.570000 39.020000 151.440000 ;
      RECT 0.000000 150.330000 40.020000 150.570000 ;
      RECT 1.000000 149.800000 40.020000 150.330000 ;
      RECT 39.290000 149.720000 40.020000 149.800000 ;
      RECT 39.290000 148.720000 40.020000 148.740000 ;
      RECT 6.560000 148.720000 37.490000 149.800000 ;
      RECT 2.530000 148.720000 4.595000 149.800000 ;
      RECT 0.000000 148.720000 0.730000 149.350000 ;
      RECT 0.000000 148.500000 40.020000 148.720000 ;
      RECT 0.000000 147.520000 39.020000 148.500000 ;
      RECT 0.000000 147.080000 40.020000 147.520000 ;
      RECT 37.490000 146.670000 40.020000 147.080000 ;
      RECT 0.000000 146.060000 2.530000 147.080000 ;
      RECT 37.490000 146.000000 39.020000 146.670000 ;
      RECT 8.560000 146.000000 35.690000 147.080000 ;
      RECT 4.330000 146.000000 6.760000 147.080000 ;
      RECT 1.000000 146.000000 2.530000 146.060000 ;
      RECT 1.000000 145.690000 39.020000 146.000000 ;
      RECT 1.000000 145.450000 40.020000 145.690000 ;
      RECT 1.000000 145.080000 39.020000 145.450000 ;
      RECT 0.000000 144.470000 39.020000 145.080000 ;
      RECT 0.000000 144.360000 40.020000 144.470000 ;
      RECT 39.290000 144.230000 40.020000 144.360000 ;
      RECT 6.560000 143.280000 37.490000 144.360000 ;
      RECT 2.530000 143.280000 4.595000 144.360000 ;
      RECT 0.000000 143.280000 0.730000 144.360000 ;
      RECT 0.000000 143.250000 39.020000 143.280000 ;
      RECT 0.000000 142.400000 40.020000 143.250000 ;
      RECT 1.000000 141.640000 39.020000 142.400000 ;
      RECT 37.490000 141.420000 39.020000 141.640000 ;
      RECT 1.000000 141.420000 2.530000 141.640000 ;
      RECT 37.490000 141.180000 40.020000 141.420000 ;
      RECT 37.490000 140.560000 39.020000 141.180000 ;
      RECT 8.560000 140.560000 35.690000 141.640000 ;
      RECT 4.330000 140.560000 6.760000 141.640000 ;
      RECT 0.000000 140.560000 2.530000 141.420000 ;
      RECT 0.000000 140.200000 39.020000 140.560000 ;
      RECT 0.000000 139.350000 40.020000 140.200000 ;
      RECT 0.000000 138.920000 39.020000 139.350000 ;
      RECT 0.000000 138.740000 0.730000 138.920000 ;
      RECT 39.290000 138.130000 40.020000 138.370000 ;
      RECT 6.560000 137.840000 37.490000 138.920000 ;
      RECT 2.530000 137.840000 4.595000 138.920000 ;
      RECT 1.000000 137.760000 39.020000 137.840000 ;
      RECT 0.000000 137.150000 39.020000 137.760000 ;
      RECT 0.000000 136.300000 40.020000 137.150000 ;
      RECT 0.000000 136.200000 39.020000 136.300000 ;
      RECT 37.490000 135.320000 39.020000 136.200000 ;
      RECT 37.490000 135.120000 40.020000 135.320000 ;
      RECT 8.560000 135.120000 35.690000 136.200000 ;
      RECT 4.330000 135.120000 6.760000 136.200000 ;
      RECT 0.000000 135.120000 2.530000 136.200000 ;
      RECT 0.000000 135.080000 40.020000 135.120000 ;
      RECT 1.000000 134.100000 39.020000 135.080000 ;
      RECT 0.000000 133.480000 40.020000 134.100000 ;
      RECT 39.290000 133.250000 40.020000 133.480000 ;
      RECT 6.560000 132.400000 37.490000 133.480000 ;
      RECT 2.530000 132.400000 4.595000 133.480000 ;
      RECT 0.000000 132.400000 0.730000 133.480000 ;
      RECT 0.000000 132.270000 39.020000 132.400000 ;
      RECT 0.000000 132.030000 40.020000 132.270000 ;
      RECT 0.000000 131.420000 39.020000 132.030000 ;
      RECT 1.000000 131.050000 39.020000 131.420000 ;
      RECT 1.000000 130.810000 40.020000 131.050000 ;
      RECT 1.000000 130.760000 39.020000 130.810000 ;
      RECT 1.000000 130.440000 2.530000 130.760000 ;
      RECT 37.490000 129.830000 39.020000 130.760000 ;
      RECT 37.490000 129.680000 40.020000 129.830000 ;
      RECT 8.560000 129.680000 35.690000 130.760000 ;
      RECT 4.330000 129.680000 6.760000 130.760000 ;
      RECT 0.000000 129.680000 2.530000 130.440000 ;
      RECT 0.000000 128.980000 40.020000 129.680000 ;
      RECT 0.000000 128.040000 39.020000 128.980000 ;
      RECT 39.290000 127.760000 40.020000 128.000000 ;
      RECT 0.000000 127.760000 0.730000 128.040000 ;
      RECT 6.560000 126.960000 37.490000 128.040000 ;
      RECT 2.530000 126.960000 4.595000 128.040000 ;
      RECT 1.000000 126.780000 39.020000 126.960000 ;
      RECT 0.000000 125.930000 40.020000 126.780000 ;
      RECT 0.000000 125.320000 39.020000 125.930000 ;
      RECT 37.490000 124.950000 39.020000 125.320000 ;
      RECT 37.490000 124.710000 40.020000 124.950000 ;
      RECT 37.490000 124.240000 39.020000 124.710000 ;
      RECT 8.560000 124.240000 35.690000 125.320000 ;
      RECT 4.330000 124.240000 6.760000 125.320000 ;
      RECT 0.000000 124.240000 2.530000 125.320000 ;
      RECT 0.000000 124.100000 39.020000 124.240000 ;
      RECT 1.000000 123.730000 39.020000 124.100000 ;
      RECT 1.000000 123.120000 40.020000 123.730000 ;
      RECT 0.000000 122.880000 40.020000 123.120000 ;
      RECT 0.000000 122.600000 39.020000 122.880000 ;
      RECT 39.290000 121.660000 40.020000 121.900000 ;
      RECT 6.560000 121.520000 37.490000 122.600000 ;
      RECT 2.530000 121.520000 4.595000 122.600000 ;
      RECT 0.000000 121.520000 0.730000 122.600000 ;
      RECT 0.000000 120.680000 39.020000 121.520000 ;
      RECT 0.000000 120.440000 40.020000 120.680000 ;
      RECT 1.000000 119.880000 40.020000 120.440000 ;
      RECT 37.490000 119.830000 40.020000 119.880000 ;
      RECT 1.000000 119.460000 2.530000 119.880000 ;
      RECT 37.490000 118.850000 39.020000 119.830000 ;
      RECT 37.490000 118.800000 40.020000 118.850000 ;
      RECT 8.560000 118.800000 35.690000 119.880000 ;
      RECT 4.330000 118.800000 6.760000 119.880000 ;
      RECT 0.000000 118.800000 2.530000 119.460000 ;
      RECT 0.000000 118.610000 40.020000 118.800000 ;
      RECT 0.000000 117.630000 39.020000 118.610000 ;
      RECT 0.000000 117.390000 40.020000 117.630000 ;
      RECT 0.000000 117.160000 39.020000 117.390000 ;
      RECT 0.000000 116.780000 0.730000 117.160000 ;
      RECT 39.290000 116.080000 40.020000 116.410000 ;
      RECT 6.560000 116.080000 37.490000 117.160000 ;
      RECT 2.530000 116.080000 4.595000 117.160000 ;
      RECT 1.000000 115.800000 40.020000 116.080000 ;
      RECT 0.000000 115.560000 40.020000 115.800000 ;
      RECT 0.000000 114.580000 39.020000 115.560000 ;
      RECT 0.000000 114.440000 40.020000 114.580000 ;
      RECT 37.490000 114.340000 40.020000 114.440000 ;
      RECT 37.490000 113.360000 39.020000 114.340000 ;
      RECT 8.560000 113.360000 35.690000 114.440000 ;
      RECT 4.330000 113.360000 6.760000 114.440000 ;
      RECT 0.000000 113.360000 2.530000 114.440000 ;
      RECT 0.000000 113.120000 40.020000 113.360000 ;
      RECT 1.000000 112.510000 40.020000 113.120000 ;
      RECT 1.000000 112.140000 39.020000 112.510000 ;
      RECT 0.000000 111.720000 39.020000 112.140000 ;
      RECT 39.290000 111.290000 40.020000 111.530000 ;
      RECT 6.560000 110.640000 37.490000 111.720000 ;
      RECT 2.530000 110.640000 4.595000 111.720000 ;
      RECT 0.000000 110.640000 0.730000 111.720000 ;
      RECT 0.000000 110.310000 39.020000 110.640000 ;
      RECT 0.000000 109.460000 40.020000 110.310000 ;
      RECT 1.000000 109.000000 39.020000 109.460000 ;
      RECT 37.490000 108.480000 39.020000 109.000000 ;
      RECT 1.000000 108.480000 2.530000 109.000000 ;
      RECT 37.490000 108.240000 40.020000 108.480000 ;
      RECT 37.490000 107.920000 39.020000 108.240000 ;
      RECT 8.560000 107.920000 35.690000 109.000000 ;
      RECT 4.330000 107.920000 6.760000 109.000000 ;
      RECT 0.000000 107.920000 2.530000 108.480000 ;
      RECT 0.000000 107.260000 39.020000 107.920000 ;
      RECT 0.000000 106.410000 40.020000 107.260000 ;
      RECT 0.000000 106.280000 39.020000 106.410000 ;
      RECT 0.000000 105.800000 0.730000 106.280000 ;
      RECT 39.290000 105.200000 40.020000 105.430000 ;
      RECT 6.560000 105.200000 37.490000 106.280000 ;
      RECT 2.530000 105.200000 4.595000 106.280000 ;
      RECT 1.000000 105.190000 40.020000 105.200000 ;
      RECT 1.000000 104.820000 39.020000 105.190000 ;
      RECT 0.000000 104.210000 39.020000 104.820000 ;
      RECT 0.000000 103.970000 40.020000 104.210000 ;
      RECT 0.000000 103.560000 39.020000 103.970000 ;
      RECT 37.490000 102.990000 39.020000 103.560000 ;
      RECT 37.490000 102.480000 40.020000 102.990000 ;
      RECT 8.560000 102.480000 35.690000 103.560000 ;
      RECT 4.330000 102.480000 6.760000 103.560000 ;
      RECT 0.000000 102.480000 2.530000 103.560000 ;
      RECT 0.000000 102.140000 40.020000 102.480000 ;
      RECT 1.000000 101.160000 39.020000 102.140000 ;
      RECT 0.000000 100.920000 40.020000 101.160000 ;
      RECT 0.000000 100.840000 39.020000 100.920000 ;
      RECT 39.290000 99.760000 40.020000 99.940000 ;
      RECT 6.560000 99.760000 37.490000 100.840000 ;
      RECT 2.530000 99.760000 4.595000 100.840000 ;
      RECT 0.000000 99.760000 0.730000 100.840000 ;
      RECT 0.000000 99.090000 40.020000 99.760000 ;
      RECT 0.000000 98.120000 39.020000 99.090000 ;
      RECT 37.490000 98.110000 39.020000 98.120000 ;
      RECT 37.490000 97.870000 40.020000 98.110000 ;
      RECT 0.000000 97.870000 2.530000 98.120000 ;
      RECT 37.490000 97.040000 39.020000 97.870000 ;
      RECT 8.560000 97.040000 35.690000 98.120000 ;
      RECT 4.330000 97.040000 6.760000 98.120000 ;
      RECT 1.000000 97.040000 2.530000 97.870000 ;
      RECT 1.000000 96.890000 39.020000 97.040000 ;
      RECT 0.000000 96.040000 40.020000 96.890000 ;
      RECT 0.000000 95.400000 39.020000 96.040000 ;
      RECT 39.290000 94.820000 40.020000 95.060000 ;
      RECT 6.560000 94.320000 37.490000 95.400000 ;
      RECT 2.530000 94.320000 4.595000 95.400000 ;
      RECT 0.000000 94.320000 0.730000 95.400000 ;
      RECT 0.000000 94.210000 39.020000 94.320000 ;
      RECT 1.000000 93.840000 39.020000 94.210000 ;
      RECT 1.000000 93.600000 40.020000 93.840000 ;
      RECT 1.000000 93.230000 39.020000 93.600000 ;
      RECT 0.000000 92.680000 39.020000 93.230000 ;
      RECT 37.490000 92.620000 39.020000 92.680000 ;
      RECT 37.490000 91.770000 40.020000 92.620000 ;
      RECT 37.490000 91.600000 39.020000 91.770000 ;
      RECT 8.560000 91.600000 35.690000 92.680000 ;
      RECT 4.330000 91.600000 6.760000 92.680000 ;
      RECT 0.000000 91.600000 2.530000 92.680000 ;
      RECT 0.000000 90.790000 39.020000 91.600000 ;
      RECT 0.000000 90.550000 40.020000 90.790000 ;
      RECT 1.000000 89.960000 39.020000 90.550000 ;
      RECT 39.290000 88.880000 40.020000 89.570000 ;
      RECT 6.560000 88.880000 37.490000 89.960000 ;
      RECT 2.530000 88.880000 4.595000 89.960000 ;
      RECT 0.000000 88.880000 0.730000 89.570000 ;
      RECT 0.000000 88.720000 40.020000 88.880000 ;
      RECT 0.000000 87.740000 39.020000 88.720000 ;
      RECT 0.000000 87.500000 40.020000 87.740000 ;
      RECT 0.000000 87.240000 39.020000 87.500000 ;
      RECT 0.000000 86.890000 2.530000 87.240000 ;
      RECT 37.490000 86.520000 39.020000 87.240000 ;
      RECT 37.490000 86.160000 40.020000 86.520000 ;
      RECT 8.560000 86.160000 35.690000 87.240000 ;
      RECT 4.330000 86.160000 6.760000 87.240000 ;
      RECT 1.000000 86.160000 2.530000 86.890000 ;
      RECT 1.000000 85.910000 40.020000 86.160000 ;
      RECT 0.000000 85.670000 40.020000 85.910000 ;
      RECT 0.000000 84.690000 39.020000 85.670000 ;
      RECT 0.000000 84.520000 40.020000 84.690000 ;
      RECT 39.290000 84.450000 40.020000 84.520000 ;
      RECT 39.290000 83.440000 40.020000 83.470000 ;
      RECT 6.560000 83.440000 37.490000 84.520000 ;
      RECT 2.530000 83.440000 4.595000 84.520000 ;
      RECT 0.000000 83.440000 0.730000 84.520000 ;
      RECT 0.000000 83.230000 40.020000 83.440000 ;
      RECT 1.000000 82.620000 40.020000 83.230000 ;
      RECT 1.000000 82.250000 39.020000 82.620000 ;
      RECT 0.000000 81.800000 39.020000 82.250000 ;
      RECT 37.490000 81.640000 39.020000 81.800000 ;
      RECT 37.490000 81.400000 40.020000 81.640000 ;
      RECT 37.490000 80.720000 39.020000 81.400000 ;
      RECT 8.560000 80.720000 35.690000 81.800000 ;
      RECT 4.330000 80.720000 6.760000 81.800000 ;
      RECT 0.000000 80.720000 2.530000 81.800000 ;
      RECT 0.000000 80.420000 39.020000 80.720000 ;
      RECT 0.000000 80.180000 40.020000 80.420000 ;
      RECT 0.000000 79.570000 39.020000 80.180000 ;
      RECT 1.000000 79.200000 39.020000 79.570000 ;
      RECT 1.000000 79.080000 40.020000 79.200000 ;
      RECT 39.290000 78.350000 40.020000 79.080000 ;
      RECT 6.560000 78.000000 37.490000 79.080000 ;
      RECT 2.530000 78.000000 4.595000 79.080000 ;
      RECT 0.000000 78.000000 0.730000 78.590000 ;
      RECT 0.000000 77.370000 39.020000 78.000000 ;
      RECT 0.000000 77.130000 40.020000 77.370000 ;
      RECT 0.000000 76.360000 39.020000 77.130000 ;
      RECT 37.490000 76.150000 39.020000 76.360000 ;
      RECT 0.000000 75.910000 2.530000 76.360000 ;
      RECT 37.490000 75.300000 40.020000 76.150000 ;
      RECT 37.490000 75.280000 39.020000 75.300000 ;
      RECT 8.560000 75.280000 35.690000 76.360000 ;
      RECT 4.330000 75.280000 6.760000 76.360000 ;
      RECT 1.000000 75.280000 2.530000 75.910000 ;
      RECT 1.000000 74.930000 39.020000 75.280000 ;
      RECT 0.000000 74.320000 39.020000 74.930000 ;
      RECT 0.000000 74.080000 40.020000 74.320000 ;
      RECT 0.000000 73.640000 39.020000 74.080000 ;
      RECT 39.290000 72.560000 40.020000 73.100000 ;
      RECT 6.560000 72.560000 37.490000 73.640000 ;
      RECT 2.530000 72.560000 4.595000 73.640000 ;
      RECT 0.000000 72.560000 0.730000 73.640000 ;
      RECT 0.000000 72.250000 40.020000 72.560000 ;
      RECT 1.000000 71.270000 39.020000 72.250000 ;
      RECT 0.000000 71.030000 40.020000 71.270000 ;
      RECT 0.000000 70.920000 39.020000 71.030000 ;
      RECT 37.490000 70.050000 39.020000 70.920000 ;
      RECT 37.490000 69.840000 40.020000 70.050000 ;
      RECT 8.560000 69.840000 35.690000 70.920000 ;
      RECT 4.330000 69.840000 6.760000 70.920000 ;
      RECT 0.000000 69.840000 2.530000 70.920000 ;
      RECT 0.000000 69.200000 40.020000 69.840000 ;
      RECT 0.000000 68.590000 39.020000 69.200000 ;
      RECT 1.000000 68.220000 39.020000 68.590000 ;
      RECT 1.000000 68.200000 40.020000 68.220000 ;
      RECT 39.290000 67.980000 40.020000 68.200000 ;
      RECT 6.560000 67.120000 37.490000 68.200000 ;
      RECT 2.530000 67.120000 4.595000 68.200000 ;
      RECT 0.000000 67.120000 0.730000 67.610000 ;
      RECT 0.000000 67.000000 39.020000 67.120000 ;
      RECT 0.000000 66.760000 40.020000 67.000000 ;
      RECT 0.000000 65.780000 39.020000 66.760000 ;
      RECT 0.000000 65.480000 40.020000 65.780000 ;
      RECT 37.490000 64.930000 40.020000 65.480000 ;
      RECT 0.000000 64.930000 2.530000 65.480000 ;
      RECT 37.490000 64.400000 39.020000 64.930000 ;
      RECT 8.560000 64.400000 35.690000 65.480000 ;
      RECT 4.330000 64.400000 6.760000 65.480000 ;
      RECT 1.000000 64.400000 2.530000 64.930000 ;
      RECT 1.000000 63.950000 39.020000 64.400000 ;
      RECT 0.000000 63.710000 40.020000 63.950000 ;
      RECT 0.000000 62.760000 39.020000 63.710000 ;
      RECT 39.290000 61.880000 40.020000 62.730000 ;
      RECT 6.560000 61.680000 37.490000 62.760000 ;
      RECT 2.530000 61.680000 4.595000 62.760000 ;
      RECT 0.000000 61.680000 0.730000 62.760000 ;
      RECT 0.000000 61.270000 39.020000 61.680000 ;
      RECT 1.000000 60.900000 39.020000 61.270000 ;
      RECT 1.000000 60.660000 40.020000 60.900000 ;
      RECT 1.000000 60.290000 39.020000 60.660000 ;
      RECT 0.000000 60.040000 39.020000 60.290000 ;
      RECT 37.490000 59.680000 39.020000 60.040000 ;
      RECT 37.490000 58.960000 40.020000 59.680000 ;
      RECT 8.560000 58.960000 35.690000 60.040000 ;
      RECT 4.330000 58.960000 6.760000 60.040000 ;
      RECT 0.000000 58.960000 2.530000 60.040000 ;
      RECT 0.000000 58.830000 40.020000 58.960000 ;
      RECT 0.000000 57.850000 39.020000 58.830000 ;
      RECT 0.000000 57.610000 40.020000 57.850000 ;
      RECT 1.000000 57.320000 39.020000 57.610000 ;
      RECT 39.290000 56.240000 40.020000 56.630000 ;
      RECT 6.560000 56.240000 37.490000 57.320000 ;
      RECT 2.530000 56.240000 4.595000 57.320000 ;
      RECT 0.000000 56.240000 0.730000 56.630000 ;
      RECT 0.000000 55.780000 40.020000 56.240000 ;
      RECT 0.000000 54.800000 39.020000 55.780000 ;
      RECT 0.000000 54.600000 40.020000 54.800000 ;
      RECT 37.490000 54.560000 40.020000 54.600000 ;
      RECT 0.000000 53.950000 2.530000 54.600000 ;
      RECT 37.490000 53.580000 39.020000 54.560000 ;
      RECT 37.490000 53.520000 40.020000 53.580000 ;
      RECT 8.560000 53.520000 35.690000 54.600000 ;
      RECT 4.330000 53.520000 6.760000 54.600000 ;
      RECT 1.000000 53.520000 2.530000 53.950000 ;
      RECT 1.000000 53.340000 40.020000 53.520000 ;
      RECT 1.000000 52.970000 39.020000 53.340000 ;
      RECT 0.000000 52.360000 39.020000 52.970000 ;
      RECT 0.000000 51.880000 40.020000 52.360000 ;
      RECT 39.290000 51.510000 40.020000 51.880000 ;
      RECT 6.560000 50.800000 37.490000 51.880000 ;
      RECT 2.530000 50.800000 4.595000 51.880000 ;
      RECT 0.000000 50.800000 0.730000 51.880000 ;
      RECT 0.000000 50.530000 39.020000 50.800000 ;
      RECT 0.000000 50.290000 40.020000 50.530000 ;
      RECT 0.000000 49.680000 39.020000 50.290000 ;
      RECT 1.000000 49.310000 39.020000 49.680000 ;
      RECT 1.000000 49.160000 40.020000 49.310000 ;
      RECT 1.000000 48.700000 2.530000 49.160000 ;
      RECT 37.490000 48.460000 40.020000 49.160000 ;
      RECT 37.490000 48.080000 39.020000 48.460000 ;
      RECT 8.560000 48.080000 35.690000 49.160000 ;
      RECT 4.330000 48.080000 6.760000 49.160000 ;
      RECT 0.000000 48.080000 2.530000 48.700000 ;
      RECT 0.000000 47.480000 39.020000 48.080000 ;
      RECT 0.000000 47.240000 40.020000 47.480000 ;
      RECT 0.000000 46.440000 39.020000 47.240000 ;
      RECT 0.000000 46.020000 0.730000 46.440000 ;
      RECT 39.290000 45.410000 40.020000 46.260000 ;
      RECT 6.560000 45.360000 37.490000 46.440000 ;
      RECT 2.530000 45.360000 4.595000 46.440000 ;
      RECT 1.000000 45.040000 39.020000 45.360000 ;
      RECT 0.000000 44.430000 39.020000 45.040000 ;
      RECT 0.000000 44.190000 40.020000 44.430000 ;
      RECT 0.000000 43.720000 39.020000 44.190000 ;
      RECT 37.490000 43.210000 39.020000 43.720000 ;
      RECT 37.490000 42.970000 40.020000 43.210000 ;
      RECT 37.490000 42.640000 39.020000 42.970000 ;
      RECT 8.560000 42.640000 35.690000 43.720000 ;
      RECT 4.330000 42.640000 6.760000 43.720000 ;
      RECT 0.000000 42.640000 2.530000 43.720000 ;
      RECT 0.000000 42.360000 39.020000 42.640000 ;
      RECT 1.000000 41.990000 39.020000 42.360000 ;
      RECT 1.000000 41.380000 40.020000 41.990000 ;
      RECT 0.000000 41.140000 40.020000 41.380000 ;
      RECT 0.000000 41.000000 39.020000 41.140000 ;
      RECT 39.290000 39.920000 40.020000 40.160000 ;
      RECT 6.560000 39.920000 37.490000 41.000000 ;
      RECT 2.530000 39.920000 4.595000 41.000000 ;
      RECT 0.000000 39.920000 0.730000 41.000000 ;
      RECT 0.000000 38.940000 39.020000 39.920000 ;
      RECT 0.000000 38.700000 40.020000 38.940000 ;
      RECT 1.000000 38.280000 40.020000 38.700000 ;
      RECT 37.490000 38.090000 40.020000 38.280000 ;
      RECT 1.000000 37.720000 2.530000 38.280000 ;
      RECT 37.490000 37.200000 39.020000 38.090000 ;
      RECT 8.560000 37.200000 35.690000 38.280000 ;
      RECT 4.330000 37.200000 6.760000 38.280000 ;
      RECT 0.000000 37.200000 2.530000 37.720000 ;
      RECT 0.000000 37.110000 39.020000 37.200000 ;
      RECT 0.000000 36.870000 40.020000 37.110000 ;
      RECT 0.000000 35.890000 39.020000 36.870000 ;
      RECT 0.000000 35.560000 40.020000 35.890000 ;
      RECT 39.290000 35.040000 40.020000 35.560000 ;
      RECT 0.000000 35.040000 0.730000 35.560000 ;
      RECT 6.560000 34.480000 37.490000 35.560000 ;
      RECT 2.530000 34.480000 4.595000 35.560000 ;
      RECT 1.000000 34.060000 39.020000 34.480000 ;
      RECT 0.000000 33.820000 40.020000 34.060000 ;
      RECT 0.000000 32.840000 39.020000 33.820000 ;
      RECT 37.490000 31.990000 40.020000 32.840000 ;
      RECT 37.490000 31.760000 39.020000 31.990000 ;
      RECT 8.560000 31.760000 35.690000 32.840000 ;
      RECT 4.330000 31.760000 6.760000 32.840000 ;
      RECT 0.000000 31.760000 2.530000 32.840000 ;
      RECT 0.000000 31.380000 39.020000 31.760000 ;
      RECT 1.000000 31.010000 39.020000 31.380000 ;
      RECT 1.000000 30.770000 40.020000 31.010000 ;
      RECT 1.000000 30.400000 39.020000 30.770000 ;
      RECT 0.000000 30.120000 39.020000 30.400000 ;
      RECT 39.290000 29.550000 40.020000 29.790000 ;
      RECT 6.560000 29.040000 37.490000 30.120000 ;
      RECT 2.530000 29.040000 4.595000 30.120000 ;
      RECT 0.000000 29.040000 0.730000 30.120000 ;
      RECT 0.000000 28.570000 39.020000 29.040000 ;
      RECT 0.000000 27.720000 40.020000 28.570000 ;
      RECT 1.000000 27.400000 39.020000 27.720000 ;
      RECT 37.490000 26.740000 39.020000 27.400000 ;
      RECT 1.000000 26.740000 2.530000 27.400000 ;
      RECT 37.490000 26.500000 40.020000 26.740000 ;
      RECT 37.490000 26.320000 39.020000 26.500000 ;
      RECT 8.560000 26.320000 35.690000 27.400000 ;
      RECT 4.330000 26.320000 6.760000 27.400000 ;
      RECT 0.000000 26.320000 2.530000 26.740000 ;
      RECT 0.000000 25.520000 39.020000 26.320000 ;
      RECT 0.000000 24.680000 40.020000 25.520000 ;
      RECT 39.290000 24.670000 40.020000 24.680000 ;
      RECT 0.000000 24.060000 0.730000 24.680000 ;
      RECT 39.290000 23.600000 40.020000 23.690000 ;
      RECT 6.560000 23.600000 37.490000 24.680000 ;
      RECT 2.530000 23.600000 4.595000 24.680000 ;
      RECT 1.000000 23.450000 40.020000 23.600000 ;
      RECT 1.000000 23.080000 39.020000 23.450000 ;
      RECT 0.000000 22.470000 39.020000 23.080000 ;
      RECT 0.000000 21.960000 40.020000 22.470000 ;
      RECT 37.490000 21.620000 40.020000 21.960000 ;
      RECT 37.490000 20.880000 39.020000 21.620000 ;
      RECT 8.560000 20.880000 35.690000 21.960000 ;
      RECT 4.330000 20.880000 6.760000 21.960000 ;
      RECT 0.000000 20.880000 2.530000 21.960000 ;
      RECT 0.000000 20.640000 39.020000 20.880000 ;
      RECT 0.000000 20.400000 40.020000 20.640000 ;
      RECT 1.000000 19.420000 39.020000 20.400000 ;
      RECT 0.000000 19.240000 40.020000 19.420000 ;
      RECT 39.290000 18.570000 40.020000 19.240000 ;
      RECT 6.560000 18.160000 37.490000 19.240000 ;
      RECT 2.530000 18.160000 4.595000 19.240000 ;
      RECT 0.000000 18.160000 0.730000 19.240000 ;
      RECT 0.000000 17.590000 39.020000 18.160000 ;
      RECT 0.000000 17.350000 40.020000 17.590000 ;
      RECT 0.000000 16.740000 39.020000 17.350000 ;
      RECT 1.000000 16.520000 39.020000 16.740000 ;
      RECT 37.490000 16.370000 39.020000 16.520000 ;
      RECT 37.490000 16.130000 40.020000 16.370000 ;
      RECT 1.000000 15.760000 2.530000 16.520000 ;
      RECT 37.490000 15.440000 39.020000 16.130000 ;
      RECT 8.560000 15.440000 35.690000 16.520000 ;
      RECT 4.330000 15.440000 6.760000 16.520000 ;
      RECT 0.000000 15.440000 2.530000 15.760000 ;
      RECT 0.000000 15.150000 39.020000 15.440000 ;
      RECT 0.000000 14.300000 40.020000 15.150000 ;
      RECT 0.000000 13.800000 39.020000 14.300000 ;
      RECT 39.290000 13.080000 40.020000 13.320000 ;
      RECT 0.000000 13.080000 0.730000 13.800000 ;
      RECT 6.560000 12.720000 37.490000 13.800000 ;
      RECT 2.530000 12.720000 4.595000 13.800000 ;
      RECT 1.000000 12.100000 39.020000 12.720000 ;
      RECT 0.000000 11.250000 40.020000 12.100000 ;
      RECT 0.000000 11.080000 39.020000 11.250000 ;
      RECT 37.490000 10.270000 39.020000 11.080000 ;
      RECT 37.490000 10.030000 40.020000 10.270000 ;
      RECT 37.490000 10.000000 39.020000 10.030000 ;
      RECT 8.560000 10.000000 35.690000 11.080000 ;
      RECT 4.330000 10.000000 6.760000 11.080000 ;
      RECT 0.000000 10.000000 2.530000 11.080000 ;
      RECT 0.000000 9.420000 39.020000 10.000000 ;
      RECT 1.000000 9.050000 39.020000 9.420000 ;
      RECT 1.000000 8.440000 40.020000 9.050000 ;
      RECT 0.000000 8.360000 40.020000 8.440000 ;
      RECT 39.290000 8.200000 40.020000 8.360000 ;
      RECT 6.560000 7.280000 37.490000 8.360000 ;
      RECT 2.530000 7.280000 4.595000 8.360000 ;
      RECT 0.000000 7.280000 0.730000 8.360000 ;
      RECT 0.000000 7.220000 39.020000 7.280000 ;
      RECT 0.000000 6.980000 40.020000 7.220000 ;
      RECT 0.000000 6.000000 39.020000 6.980000 ;
      RECT 0.000000 5.760000 40.020000 6.000000 ;
      RECT 1.000000 5.640000 39.020000 5.760000 ;
      RECT 37.490000 4.780000 39.020000 5.640000 ;
      RECT 1.000000 4.780000 2.530000 5.640000 ;
      RECT 37.490000 4.560000 40.020000 4.780000 ;
      RECT 8.560000 4.560000 35.690000 5.640000 ;
      RECT 4.330000 4.560000 6.760000 5.640000 ;
      RECT 0.000000 4.560000 2.530000 4.780000 ;
      RECT 0.000000 4.350000 40.020000 4.560000 ;
      RECT 0.000000 0.000000 40.020000 0.750000 ;
    LAYER met4 ;
      RECT 4.330000 198.320000 35.690000 200.260000 ;
      RECT 6.560000 196.520000 35.690000 198.320000 ;
      RECT 4.330000 193.320000 4.760000 198.320000 ;
      RECT 4.330000 192.240000 4.595000 193.320000 ;
      RECT 4.330000 187.880000 4.760000 192.240000 ;
      RECT 4.330000 186.800000 4.595000 187.880000 ;
      RECT 4.330000 182.440000 4.760000 186.800000 ;
      RECT 4.330000 181.360000 4.595000 182.440000 ;
      RECT 4.330000 177.000000 4.760000 181.360000 ;
      RECT 4.330000 175.920000 4.595000 177.000000 ;
      RECT 4.330000 171.560000 4.760000 175.920000 ;
      RECT 4.330000 170.480000 4.595000 171.560000 ;
      RECT 4.330000 166.120000 4.760000 170.480000 ;
      RECT 4.330000 165.040000 4.595000 166.120000 ;
      RECT 4.330000 160.680000 4.760000 165.040000 ;
      RECT 4.330000 159.600000 4.595000 160.680000 ;
      RECT 4.330000 155.240000 4.760000 159.600000 ;
      RECT 4.330000 154.160000 4.595000 155.240000 ;
      RECT 4.330000 149.800000 4.760000 154.160000 ;
      RECT 4.330000 148.720000 4.595000 149.800000 ;
      RECT 4.330000 144.360000 4.760000 148.720000 ;
      RECT 4.330000 143.280000 4.595000 144.360000 ;
      RECT 4.330000 138.920000 4.760000 143.280000 ;
      RECT 4.330000 137.840000 4.595000 138.920000 ;
      RECT 4.330000 133.480000 4.760000 137.840000 ;
      RECT 4.330000 132.400000 4.595000 133.480000 ;
      RECT 4.330000 128.040000 4.760000 132.400000 ;
      RECT 4.330000 126.960000 4.595000 128.040000 ;
      RECT 4.330000 122.600000 4.760000 126.960000 ;
      RECT 4.330000 121.520000 4.595000 122.600000 ;
      RECT 4.330000 117.160000 4.760000 121.520000 ;
      RECT 4.330000 116.080000 4.595000 117.160000 ;
      RECT 4.330000 111.720000 4.760000 116.080000 ;
      RECT 4.330000 110.640000 4.595000 111.720000 ;
      RECT 4.330000 106.280000 4.760000 110.640000 ;
      RECT 4.330000 105.200000 4.595000 106.280000 ;
      RECT 4.330000 100.840000 4.760000 105.200000 ;
      RECT 4.330000 99.760000 4.595000 100.840000 ;
      RECT 4.330000 95.400000 4.760000 99.760000 ;
      RECT 4.330000 94.320000 4.595000 95.400000 ;
      RECT 4.330000 89.960000 4.760000 94.320000 ;
      RECT 4.330000 88.880000 4.595000 89.960000 ;
      RECT 4.330000 84.520000 4.760000 88.880000 ;
      RECT 4.330000 83.440000 4.595000 84.520000 ;
      RECT 4.330000 79.080000 4.760000 83.440000 ;
      RECT 4.330000 78.000000 4.595000 79.080000 ;
      RECT 4.330000 73.640000 4.760000 78.000000 ;
      RECT 4.330000 72.560000 4.595000 73.640000 ;
      RECT 4.330000 68.200000 4.760000 72.560000 ;
      RECT 4.330000 67.120000 4.595000 68.200000 ;
      RECT 4.330000 62.760000 4.760000 67.120000 ;
      RECT 4.330000 61.680000 4.595000 62.760000 ;
      RECT 4.330000 57.320000 4.760000 61.680000 ;
      RECT 4.330000 56.240000 4.595000 57.320000 ;
      RECT 4.330000 51.880000 4.760000 56.240000 ;
      RECT 4.330000 50.800000 4.595000 51.880000 ;
      RECT 4.330000 46.440000 4.760000 50.800000 ;
      RECT 4.330000 45.360000 4.595000 46.440000 ;
      RECT 4.330000 41.000000 4.760000 45.360000 ;
      RECT 4.330000 39.920000 4.595000 41.000000 ;
      RECT 4.330000 35.560000 4.760000 39.920000 ;
      RECT 4.330000 34.480000 4.595000 35.560000 ;
      RECT 4.330000 30.120000 4.760000 34.480000 ;
      RECT 4.330000 29.040000 4.595000 30.120000 ;
      RECT 4.330000 24.680000 4.760000 29.040000 ;
      RECT 4.330000 23.600000 4.595000 24.680000 ;
      RECT 4.330000 19.240000 4.760000 23.600000 ;
      RECT 4.330000 18.160000 4.595000 19.240000 ;
      RECT 4.330000 13.800000 4.760000 18.160000 ;
      RECT 4.330000 12.720000 4.595000 13.800000 ;
      RECT 4.330000 8.360000 4.760000 12.720000 ;
      RECT 4.330000 7.280000 4.595000 8.360000 ;
      RECT 8.560000 2.550000 35.690000 196.520000 ;
      RECT 6.560000 2.550000 6.760000 196.520000 ;
      RECT 6.560000 0.750000 35.690000 2.550000 ;
      RECT 4.330000 0.750000 4.760000 7.280000 ;
      RECT 39.290000 0.000000 40.020000 200.260000 ;
      RECT 4.330000 0.000000 35.690000 0.750000 ;
      RECT 0.000000 0.000000 0.730000 200.260000 ;
  END
END W_CPU_IO

END LIBRARY
