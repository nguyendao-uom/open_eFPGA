##
## LEF for PtnCells ;
## created by Innovus v19.11-s128_1 on Mon Dec  6 20:55:28 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RegFile
  CLASS BLOCK ;
  SIZE 200.100000 BY 200.260000 ;
  FOREIGN RegFile 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.251 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 9.240000 199.560000 9.620000 200.260000 ;
    END
  END N1BEG[3]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.5854 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.701 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 7.860000 199.560000 8.240000 200.260000 ;
    END
  END N1BEG[2]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.837 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 6.480000 199.560000 6.860000 200.260000 ;
    END
  END N1BEG[1]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8897 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.0048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.496 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 199.560000 5.480000 200.260000 ;
    END
  END N1BEG[0]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.791 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.729 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 21.660000 199.560000 22.040000 200.260000 ;
    END
  END N2BEG[7]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8906 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.345 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 20.280000 199.560000 20.660000 200.260000 ;
    END
  END N2BEG[6]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6218 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.001 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 18.440000 199.560000 18.820000 200.260000 ;
    END
  END N2BEG[5]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1766 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.775 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 17.060000 199.560000 17.440000 200.260000 ;
    END
  END N2BEG[4]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.2266 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.025 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 15.680000 199.560000 16.060000 200.260000 ;
    END
  END N2BEG[3]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3626 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.587 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 13.840000 199.560000 14.220000 200.260000 ;
    END
  END N2BEG[2]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.527 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 12.460000 199.560000 12.840000 200.260000 ;
    END
  END N2BEG[1]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6526 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.155 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 11.080000 199.560000 11.460000 200.260000 ;
    END
  END N2BEG[0]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9978 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.763 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 34.080000 199.560000 34.460000 200.260000 ;
    END
  END N2BEGb[7]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.251 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 32.240000 199.560000 32.620000 200.260000 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.143 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 30.860000 199.560000 31.240000 200.260000 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5122 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.453 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 29.480000 199.560000 29.860000 200.260000 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.971 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.747 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 27.640000 199.560000 28.020000 200.260000 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0362 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.073 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 26.260000 199.560000 26.640000 200.260000 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.751 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 24.880000 199.560000 25.260000 200.260000 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8626 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.205 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 23.040000 199.560000 23.420000 200.260000 ;
    END
  END N2BEGb[0]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.168 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 58.460000 199.560000 58.840000 200.260000 ;
    END
  END N4BEG[15]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0814 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.299 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 56.620000 199.560000 57.000000 200.260000 ;
    END
  END N4BEG[14]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9145 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.058 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.4298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 88.096 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 55.240000 199.560000 55.620000 200.260000 ;
    END
  END N4BEG[13]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.5514 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.531 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 53.860000 199.560000 54.240000 200.260000 ;
    END
  END N4BEG[12]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.6158 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.853 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 52.480000 199.560000 52.860000 200.260000 ;
    END
  END N4BEG[11]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.5674 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.611 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 50.640000 199.560000 51.020000 200.260000 ;
    END
  END N4BEG[10]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.885 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.317 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 49.260000 199.560000 49.640000 200.260000 ;
    END
  END N4BEG[9]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9011 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.3445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.205 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.8768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 47.880000 199.560000 48.260000 200.260000 ;
    END
  END N4BEG[8]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4021 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.6368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 46.040000 199.560000 46.420000 200.260000 ;
    END
  END N4BEG[7]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.636 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.954 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 44.660000 199.560000 45.040000 200.260000 ;
    END
  END N4BEG[6]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.961 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.461 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 43.280000 199.560000 43.660000 200.260000 ;
    END
  END N4BEG[5]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.9695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.9488 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.864 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 41.440000 199.560000 41.820000 200.260000 ;
    END
  END N4BEG[4]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0814 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.299 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 40.060000 199.560000 40.440000 200.260000 ;
    END
  END N4BEG[3]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6831 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.3038 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.424 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 38.680000 199.560000 39.060000 200.260000 ;
    END
  END N4BEG[2]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.235 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.949 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 36.840000 199.560000 37.220000 200.260000 ;
    END
  END N4BEG[1]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2982 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.265 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 35.460000 199.560000 35.840000 200.260000 ;
    END
  END N4BEG[0]
  PIN NN4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6314 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.931 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 82.840000 199.560000 83.220000 200.260000 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9366 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.457 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 81.460000 199.560000 81.840000 200.260000 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.679 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.169 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 79.620000 199.560000 80.000000 200.260000 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.085 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 78.240000 199.560000 78.620000 200.260000 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.813 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 76.860000 199.560000 77.240000 200.260000 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.679 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.169 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 75.020000 199.560000 75.400000 200.260000 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.203 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.789 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 73.640000 199.560000 74.020000 200.260000 ;
    END
  END NN4BEG[9]
  PIN NN4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.088 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.332 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 72.260000 199.560000 72.640000 200.260000 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.733 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 70.420000 199.560000 70.800000 200.260000 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 69.040000 199.560000 69.420000 200.260000 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4006 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.895 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 67.660000 199.560000 68.040000 200.260000 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0334 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.059 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 65.820000 199.560000 66.200000 200.260000 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0194 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.989 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 64.440000 199.560000 64.820000 200.260000 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4622 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.203 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 63.060000 199.560000 63.440000 200.260000 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2982 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.265 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 61.220000 199.560000 61.600000 200.260000 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.739 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 59.840000 199.560000 60.220000 200.260000 ;
    END
  END NN4BEG[0]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5109 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.3935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.0748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.536 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3095 LAYER met4  ;
    ANTENNAMAXAREACAR 57.2469 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 283.484 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.998471 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 9.240000 0.000000 9.620000 0.700000 ;
    END
  END N1END[3]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1188 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.325 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.5226 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.6321 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.481 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.032 LAYER met3  ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 77.1516 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 398.588 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.5133 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 180.144 LAYER met4  ;
    ANTENNAGATEAREA 1.3095 LAYER met4  ;
    ANTENNAMAXAREACAR 102.744 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 536.155 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 7.860000 0.000000 8.240000 0.700000 ;
    END
  END N1END[2]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.9242 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 108.591 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met2  ;
    ANTENNAMAXAREACAR 56.6393 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 272.608 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.943 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.296 LAYER met3  ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 83.2792 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 416.156 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.6548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.168 LAYER met4  ;
    ANTENNAGATEAREA 1.3095 LAYER met4  ;
    ANTENNAMAXAREACAR 93.7067 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 473.558 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 6.480000 0.000000 6.860000 0.700000 ;
    END
  END N1END[1]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7175 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.17 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.04 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 47.7483 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 256.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3095 LAYER met4  ;
    ANTENNAMAXAREACAR 73.303 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 376.377 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 0.000000 5.480000 0.700000 ;
    END
  END N1END[0]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0518 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.819 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.51985 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.3972 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 292 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7335 LAYER met4  ;
    ANTENNAMAXAREACAR 97.604 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 505.965 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 21.660000 0.000000 22.040000 0.700000 ;
    END
  END N2MID[7]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3412 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.256 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.7689 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 1.7388 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 74.7009 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 403.104 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3133 LAYER met4  ;
    ANTENNAMAXAREACAR 56.4401 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 286.55 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.831217 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 20.280000 0.000000 20.660000 0.700000 ;
    END
  END N2MID[6]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6728 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 53.095 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 55.5552 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 273.962 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.16 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.32 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 71.6366 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 362.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.816 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 38.704 LAYER met4  ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 79.824 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 408.596 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 18.440000 0.000000 18.820000 0.700000 ;
    END
  END N2MID[5]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.0767 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.4165 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met2  ;
    ANTENNAMAXAREACAR 32.6277 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 151.91 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.548637 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAGATEAREA 0.477 LAYER met3  ;
    ANTENNAMAXAREACAR 33.1915 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 155.751 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.632495 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 23.4558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 125.568 LAYER met4  ;
    ANTENNAGATEAREA 0.6735 LAYER met4  ;
    ANTENNAMAXAREACAR 68.0182 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 342.191 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 17.060000 0.000000 17.440000 0.700000 ;
    END
  END N2MID[4]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5411 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.4575 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 31.6789 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 154.26 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.827 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.544 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 61.3328 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 314.789 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.8976 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.728 LAYER met4  ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 66.0146 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 340.888 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 15.680000 0.000000 16.060000 0.700000 ;
    END
  END N2MID[3]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7785 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.7315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.1554 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 98.24 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met4  ;
    ANTENNAMAXAREACAR 68.3046 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 355.331 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.872265 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 13.840000 0.000000 14.220000 0.700000 ;
    END
  END N2MID[2]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.484 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.151 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 36.4132 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 177.824 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.4858 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125.728 LAYER met3  ;
    ANTENNAGATEAREA 0.7995 LAYER met3  ;
    ANTENNAMAXAREACAR 65.7888 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 335.083 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 12.460000 0.000000 12.840000 0.700000 ;
    END
  END N2MID[1]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.1035 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.8945 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4815 LAYER met2  ;
    ANTENNAMAXAREACAR 43.187 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 205.673 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.547854 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.24052 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.752 LAYER met3  ;
    ANTENNAGATEAREA 0.6405 LAYER met3  ;
    ANTENNAMAXAREACAR 52.9303 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 258.369 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 11.080000 0.000000 11.460000 0.700000 ;
    END
  END N2MID[0]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.6756 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.431 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0707 LAYER met2  ;
    ANTENNAMAXAREACAR 21.2922 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 87.4321 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.360629 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.7008 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.208 LAYER met3  ;
    ANTENNAGATEAREA 1.3887 LAYER met3  ;
    ANTENNAMAXAREACAR 34.7587 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 159.592 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.449057 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 34.080000 0.000000 34.460000 0.700000 ;
    END
  END N2END[7]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2671 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0565 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 10.8496 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.4762 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.696 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 11.4026 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 39.3777 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.2357 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 201.408 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 56.9381 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 288.37 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.952201 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 32.240000 0.000000 32.620000 0.700000 ;
    END
  END N2END[6]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.2647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.5925 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met2  ;
    ANTENNAMAXAREACAR 20.2642 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 92.0606 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.376412 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.9879 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.712 LAYER met3  ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 24.6384 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 115.875 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.618717 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.4258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.408 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 45.5383 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 225.653 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.632495 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 30.860000 0.000000 31.240000 0.700000 ;
    END
  END N2END[5]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.2518 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.581 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met2  ;
    ANTENNAMAXAREACAR 14.9701 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 65.4253 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.394025 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 29.480000 0.000000 29.860000 0.700000 ;
    END
  END N2END[4]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6251 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7385 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 7.83138 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.5406 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 8.45008 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 24.755 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 61.9266 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 333.088 LAYER met4  ;
    ANTENNAGATEAREA 1.7067 LAYER met4  ;
    ANTENNAMAXAREACAR 73.2374 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 374.375 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 27.640000 0.000000 28.020000 0.700000 ;
    END
  END N2END[3]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4391 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9265 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 7.96273 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.3135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.849 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.328 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 12.2162 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 45.0725 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.7926 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 101.168 LAYER met4  ;
    ANTENNAGATEAREA 1.7067 LAYER met4  ;
    ANTENNAMAXAREACAR 47.9597 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 244.497 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.666038 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 26.260000 0.000000 26.640000 0.700000 ;
    END
  END N2END[2]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.6567 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.8865 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 16.2038 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 62.0462 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.328502 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.056 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.432 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 20.9335 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 88.3448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.42052 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.0666 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.648 LAYER met4  ;
    ANTENNAGATEAREA 1.7067 LAYER met4  ;
    ANTENNAMAXAREACAR 32.1897 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 160.564 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 24.880000 0.000000 25.260000 0.700000 ;
    END
  END N2END[1]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2263 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8625 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 7.4732 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.8659 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.047 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.384 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 32.8861 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 155.475 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.574 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 255.6 LAYER met4  ;
    ANTENNAGATEAREA 1.7067 LAYER met4  ;
    ANTENNAMAXAREACAR 61.5975 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 312.945 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 23.040000 0.000000 23.420000 0.700000 ;
    END
  END N2END[0]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.7529 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.6565 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 61.0519 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 302.265 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 58.460000 0.000000 58.840000 0.700000 ;
    END
  END N4END[15]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3231 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.4545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.04148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.5316 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.776 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 33.1934 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 176.041 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 56.620000 0.000000 57.000000 0.700000 ;
    END
  END N4END[14]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.8522 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.035 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 51.6519 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 254.237 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 55.240000 0.000000 55.620000 0.700000 ;
    END
  END N4END[13]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0419 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.7466 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 138.256 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 54.25 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 273.278 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.19033 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 53.860000 0.000000 54.240000 0.700000 ;
    END
  END N4END[12]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.0608 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.078 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 52.8941 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 260.532 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 52.480000 0.000000 52.860000 0.700000 ;
    END
  END N4END[11]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6138 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.843 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 55.5277 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 273.616 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 50.640000 0.000000 51.020000 0.700000 ;
    END
  END N4END[10]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.2466 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.007 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 59.057 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 291.346 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 49.260000 0.000000 49.640000 0.700000 ;
    END
  END N4END[9]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.6402 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.093 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 60.7323 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 300.323 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 47.880000 0.000000 48.260000 0.700000 ;
    END
  END N4END[8]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4651 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.9415 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 160.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 60.053 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 301.907 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 46.040000 0.000000 46.420000 0.700000 ;
    END
  END N4END[7]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.6381 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.0825 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 61.3771 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 303.547 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 44.660000 0.000000 45.040000 0.700000 ;
    END
  END N4END[6]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.8723 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.2535 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 56.5705 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 279.858 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 43.280000 0.000000 43.660000 0.700000 ;
    END
  END N4END[5]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.0686 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 60.235 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 62.6585 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 310.298 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 41.440000 0.000000 41.820000 0.700000 ;
    END
  END N4END[4]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5699 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5705 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 13.761 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 50.0334 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.551 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.072 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 26.5307 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 119.212 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.2842 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 270.064 LAYER met4  ;
    ANTENNAGATEAREA 1.2897 LAYER met4  ;
    ANTENNAMAXAREACAR 119.307 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 613.544 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.85635 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 40.060000 0.000000 40.440000 0.700000 ;
    END
  END N4END[3]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5035 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2485 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 8.40718 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.5358 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 10.9147 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 37.9825 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.8304 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 149.84 LAYER met4  ;
    ANTENNAGATEAREA 1.3557 LAYER met4  ;
    ANTENNAMAXAREACAR 85.2727 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 442.206 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.80021 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 38.680000 0.000000 39.060000 0.700000 ;
    END
  END N4END[2]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 18.8808 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 93.555 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1967 LAYER met2  ;
    ANTENNAMAXAREACAR 41.1032 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 197.728 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.798505 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.446 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.512 LAYER met3  ;
    ANTENNAGATEAREA 1.1967 LAYER met3  ;
    ANTENNAMAXAREACAR 43.1471 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 209.019 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.83193 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.936 LAYER met4  ;
    ANTENNAGATEAREA 1.3557 LAYER met4  ;
    ANTENNAMAXAREACAR 44.1797 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 214.873 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.83193 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 36.840000 0.000000 37.220000 0.700000 ;
    END
  END N4END[1]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.8318 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 82.901 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3557 LAYER met2  ;
    ANTENNAMAXAREACAR 29.9061 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 138.102 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 35.460000 0.000000 35.840000 0.700000 ;
    END
  END N4END[0]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.4953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 57.3685 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 59.741 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 295.71 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 82.840000 0.000000 83.220000 0.700000 ;
    END
  END NN4END[15]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.8866 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.325 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 63.2972 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 313.148 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 81.460000 0.000000 81.840000 0.700000 ;
    END
  END NN4END[14]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.4786 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 142.16 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 66.533 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 336.02 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07583 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 79.620000 0.000000 80.000000 0.700000 ;
    END
  END NN4END[13]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.257 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.177 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 54.199 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 267.656 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 78.240000 0.000000 78.620000 0.700000 ;
    END
  END NN4END[12]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1018 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 60.165 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 69.2443 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.682 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 76.860000 0.000000 77.240000 0.700000 ;
    END
  END NN4END[11]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.7962 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 68.873 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.0341 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 361.748 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 75.020000 0.000000 75.400000 0.700000 ;
    END
  END NN4END[10]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.9058 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 64.421 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 66.9191 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 331.6 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 73.640000 0.000000 74.020000 0.700000 ;
    END
  END NN4END[9]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.4607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.1955 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 56.3043 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 278.183 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 72.260000 0.000000 72.640000 0.700000 ;
    END
  END NN4END[8]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.8582 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 64.183 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 67.8687 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 335.921 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 70.420000 0.000000 70.800000 0.700000 ;
    END
  END NN4END[7]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.3182 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.483 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 58.8397 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 291.204 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 69.040000 0.000000 69.420000 0.700000 ;
    END
  END NN4END[6]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.5114 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 57.449 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 60.4046 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 298.684 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 67.660000 0.000000 68.040000 0.700000 ;
    END
  END NN4END[5]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.9882 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.833 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 53.3272 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 263.214 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 65.820000 0.000000 66.200000 0.700000 ;
    END
  END NN4END[4]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1103 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.0465 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 11.4657 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.348 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.390645 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2489 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.656 LAYER met3  ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 11.8849 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 41.1373 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.458019 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.7558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 223.168 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 92.8169 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 484.241 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700629 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 64.440000 0.000000 64.820000 0.700000 ;
    END
  END NN4END[3]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.7811 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.6365 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 23.7373 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 100.186 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.96 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 27.8321 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 123.099 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.3208 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 108.848 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 53.0834 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 267.105 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.632495 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 63.060000 0.000000 63.440000 0.700000 ;
    END
  END NN4END[2]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.1405 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 11.2774 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.5696 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.328502 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 11.864 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 41.7288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.42052 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.6764 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 265.872 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 78.0826 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 409.132 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 61.220000 0.000000 61.600000 0.700000 ;
    END
  END NN4END[1]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9877 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5515 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 29.1999 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 127.143 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 30.755 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 136.51 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 1.3041 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 54.1218 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 290.992 LAYER met4  ;
    ANTENNAGATEAREA 1.8351 LAYER met4  ;
    ANTENNAMAXAREACAR 60.2476 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 295.08 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 59.840000 0.000000 60.220000 0.700000 ;
    END
  END NN4END[0]
  PIN E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 80.720000 200.100000 81.100000 ;
    END
  END E1BEG[3]
  PIN E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.4804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.224 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 79.500000 200.100000 79.880000 ;
    END
  END E1BEG[2]
  PIN E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 77.670000 200.100000 78.050000 ;
    END
  END E1BEG[1]
  PIN E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.0786 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 76.450000 200.100000 76.830000 ;
    END
  END E1BEG[0]
  PIN E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.9024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 116.808 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 92.920000 200.100000 93.300000 ;
    END
  END E2BEG[7]
  PIN E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 91.090000 200.100000 91.470000 ;
    END
  END E2BEG[6]
  PIN E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.544 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 89.870000 200.100000 90.250000 ;
    END
  END E2BEG[5]
  PIN E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 88.040000 200.100000 88.420000 ;
    END
  END E2BEG[4]
  PIN E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 86.820000 200.100000 87.200000 ;
    END
  END E2BEG[3]
  PIN E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.656 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 84.990000 200.100000 85.370000 ;
    END
  END E2BEG[2]
  PIN E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.1264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.336 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 83.770000 200.100000 84.150000 ;
    END
  END E2BEG[1]
  PIN E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.4414 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.016 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 81.940000 200.100000 82.320000 ;
    END
  END E2BEG[0]
  PIN E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 104.510000 200.100000 104.890000 ;
    END
  END E2BEGb[7]
  PIN E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 103.290000 200.100000 103.670000 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 101.460000 200.100000 101.840000 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 100.240000 200.100000 100.620000 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 98.410000 200.100000 98.790000 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 97.190000 200.100000 97.570000 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.712 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 95.360000 200.100000 95.740000 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 94.140000 200.100000 94.520000 ;
    END
  END E2BEGb[0]
  PIN EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 128.300000 200.100000 128.680000 ;
    END
  END EE4BEG[15]
  PIN EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 127.080000 200.100000 127.460000 ;
    END
  END EE4BEG[14]
  PIN EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.1484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 125.250000 200.100000 125.630000 ;
    END
  END EE4BEG[13]
  PIN EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.896 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 124.030000 200.100000 124.410000 ;
    END
  END EE4BEG[12]
  PIN EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 122.200000 200.100000 122.580000 ;
    END
  END EE4BEG[11]
  PIN EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 120.980000 200.100000 121.360000 ;
    END
  END EE4BEG[10]
  PIN EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.1824 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.968 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 119.150000 200.100000 119.530000 ;
    END
  END EE4BEG[9]
  PIN EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.8164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.016 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 117.930000 200.100000 118.310000 ;
    END
  END EE4BEG[8]
  PIN EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 116.710000 200.100000 117.090000 ;
    END
  END EE4BEG[7]
  PIN EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 114.880000 200.100000 115.260000 ;
    END
  END EE4BEG[6]
  PIN EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 113.660000 200.100000 114.040000 ;
    END
  END EE4BEG[5]
  PIN EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 111.830000 200.100000 112.210000 ;
    END
  END EE4BEG[4]
  PIN EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.3504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 110.610000 200.100000 110.990000 ;
    END
  END EE4BEG[3]
  PIN EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8954 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.104 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 108.780000 200.100000 109.160000 ;
    END
  END EE4BEG[2]
  PIN EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.6784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 107.560000 200.100000 107.940000 ;
    END
  END EE4BEG[1]
  PIN EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 105.730000 200.100000 106.110000 ;
    END
  END EE4BEG[0]
  PIN E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.6514 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.136 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 145.990000 200.100000 146.370000 ;
    END
  END E6BEG[11]
  PIN E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4186 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.3778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 45.152 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 144.770000 200.100000 145.150000 ;
    END
  END E6BEG[10]
  PIN E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.0734 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.72 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 143.550000 200.100000 143.930000 ;
    END
  END E6BEG[9]
  PIN E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 141.720000 200.100000 142.100000 ;
    END
  END E6BEG[8]
  PIN E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 140.500000 200.100000 140.880000 ;
    END
  END E6BEG[7]
  PIN E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7634 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 138.670000 200.100000 139.050000 ;
    END
  END E6BEG[6]
  PIN E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 137.450000 200.100000 137.830000 ;
    END
  END E6BEG[5]
  PIN E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 135.620000 200.100000 136.000000 ;
    END
  END E6BEG[4]
  PIN E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 134.400000 200.100000 134.780000 ;
    END
  END E6BEG[3]
  PIN E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5514 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.936 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 132.570000 200.100000 132.950000 ;
    END
  END E6BEG[2]
  PIN E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.4024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.808 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 131.350000 200.100000 131.730000 ;
    END
  END E6BEG[1]
  PIN E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 130.130000 200.100000 130.510000 ;
    END
  END E6BEG[0]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.3436 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.44 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1505 LAYER met3  ;
    ANTENNAMAXAREACAR 47.4053 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 235.61 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 80.720000 0.700000 81.100000 ;
    END
  END E1END[3]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 59.6051 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 313.639 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 42.6006 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 228.6 LAYER met4  ;
    ANTENNAGATEAREA 1.1505 LAYER met4  ;
    ANTENNAMAXAREACAR 96.633 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 512.335 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 79.500000 0.700000 79.880000 ;
    END
  END E1END[2]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 26.6783 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 128.698 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.2195 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.3802 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 62.096 LAYER met4  ;
    ANTENNAGATEAREA 1.1505 LAYER met4  ;
    ANTENNAMAXAREACAR 72.0407 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 362.493 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.2195 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 77.670000 0.700000 78.050000 ;
    END
  END E1END[1]
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.5874 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.128 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1505 LAYER met3  ;
    ANTENNAMAXAREACAR 40.8607 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 202.263 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.641057 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 76.450000 0.700000 76.830000 ;
    END
  END E1END[0]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.3226 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 129.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.8496 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.472 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7335 LAYER met4  ;
    ANTENNAMAXAREACAR 50.2878 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 256.894 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.904061 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 92.920000 0.700000 93.300000 ;
    END
  END E2MID[7]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7136 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 25.0692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 135.584 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6585 LAYER met4  ;
    ANTENNAMAXAREACAR 96.1347 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 499.271 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.09862 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 91.090000 0.700000 91.470000 ;
    END
  END E2MID[6]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.9167 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 175.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.6938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.504 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.762 LAYER met4  ;
    ANTENNAMAXAREACAR 24.5735 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 118.378 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.691495 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 89.870000 0.700000 90.250000 ;
    END
  END E2MID[5]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6836 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.8548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 63.696 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.603 LAYER met4  ;
    ANTENNAMAXAREACAR 100.586 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 517.906 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.791732 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 88.040000 0.700000 88.420000 ;
    END
  END E2MID[4]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.6446 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 110.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.3234 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.136 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.762 LAYER met4  ;
    ANTENNAMAXAREACAR 57.5721 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 298.023 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 86.820000 0.700000 87.200000 ;
    END
  END E2MID[3]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.2876 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 140.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.603 LAYER met4  ;
    ANTENNAMAXAREACAR 16.7657 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 74.5516 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.540606 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 84.990000 0.700000 85.370000 ;
    END
  END E2MID[2]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.5356 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.051 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 130.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.729 LAYER met4  ;
    ANTENNAMAXAREACAR 136.066 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 707.02 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.67778 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 83.770000 0.700000 84.150000 ;
    END
  END E2MID[1]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8936 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.2652 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 131.296 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.57 LAYER met4  ;
    ANTENNAMAXAREACAR 114.45 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 588.426 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.36032 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 81.940000 0.700000 82.320000 ;
    END
  END E2MID[0]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.0504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.064 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0707 LAYER met3  ;
    ANTENNAMAXAREACAR 38.073 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 189.279 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.576856 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.1014 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.952 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 40.3063 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 202.206 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.576856 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 104.510000 0.700000 104.890000 ;
    END
  END E2END[7]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6596 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.4182 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 68.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 62.9393 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 323.355 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.97421 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 103.290000 0.700000 103.670000 ;
    END
  END E2END[6]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.6351 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.848 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met3  ;
    ANTENNAMAXAREACAR 36.3863 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 174.197 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 101.460000 0.700000 101.840000 ;
    END
  END E2END[5]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.6028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.352 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met3  ;
    ANTENNAMAXAREACAR 17.0023 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 67.0086 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.548637 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 100.240000 0.700000 100.620000 ;
    END
  END E2END[4]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.3551 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.488 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7997 LAYER met3  ;
    ANTENNAMAXAREACAR 33.2896 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 163.279 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.571064 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 98.410000 0.700000 98.790000 ;
    END
  END E2END[3]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.4498 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.856 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 18.7349 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 89.2318 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.642217 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.3746 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.272 LAYER met4  ;
    ANTENNAGATEAREA 1.7997 LAYER met4  ;
    ANTENNAMAXAREACAR 43.1865 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 218.608 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.771222 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 97.190000 0.700000 97.570000 ;
    END
  END E2END[2]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.3642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.408 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met3  ;
    ANTENNAMAXAREACAR 34.8696 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 169.106 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.648218 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 95.360000 0.700000 95.740000 ;
    END
  END E2END[1]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4336 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.7012 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 96.288 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 60.3373 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 313.082 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.97421 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 94.140000 0.700000 94.520000 ;
    END
  END E2END[0]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 41.9416 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 223.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.8106 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.264 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 48.8992 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 251.627 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 128.300000 0.700000 128.680000 ;
    END
  END EE4END[15]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.633 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.728 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 84.05 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 452.468 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 127.080000 0.700000 127.460000 ;
    END
  END EE4END[14]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 27.7722 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 125.675 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 125.250000 0.700000 125.630000 ;
    END
  END EE4END[13]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0434 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.9018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 87.632 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9954 LAYER met4  ;
    ANTENNAMAXAREACAR 52.0239 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 263.488 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.693294 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 124.030000 0.700000 124.410000 ;
    END
  END EE4END[12]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.257 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 92.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.8386 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 39.0154 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 210.768 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 122.200000 0.700000 122.580000 ;
    END
  END EE4END[11]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.1526 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.6712 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.128 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 45.423 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 245.302 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 120.980000 0.700000 121.360000 ;
    END
  END EE4END[10]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2854 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.984 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.0194 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 262.848 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 86.0388 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 453.303 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.324944 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 119.150000 0.700000 119.530000 ;
    END
  END EE4END[9]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.0416 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.8203 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 256.448 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 89.1347 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 456.29 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 117.930000 0.700000 118.310000 ;
    END
  END EE4END[8]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.811 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 116.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.4032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 103.669 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 557.19 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 116.710000 0.700000 117.090000 ;
    END
  END EE4END[7]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.6756 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 44.1921 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 230.553 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 114.880000 0.700000 115.260000 ;
    END
  END EE4END[6]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.71295 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.1642 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 269.424 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 109.556 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 570.6 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.729187 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 113.660000 0.700000 114.040000 ;
    END
  END EE4END[5]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5874 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.5028 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 275.152 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 98.4373 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 507.81 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.550615 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 111.830000 0.700000 112.210000 ;
    END
  END EE4END[4]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.1548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.296 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 24.9259 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 108.256 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.376412 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 110.610000 0.700000 110.990000 ;
    END
  END EE4END[3]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.8974 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.248 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 43.1226 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 208.014 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.1318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER met4  ;
    ANTENNAGATEAREA 0.7527 LAYER met4  ;
    ANTENNAMAXAREACAR 45.9548 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 223.744 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 108.780000 0.700000 109.160000 ;
    END
  END EE4END[2]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 20.2817 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 92.7122 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.517922 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 107.560000 0.700000 107.940000 ;
    END
  END EE4END[1]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 26.3731 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 113.208 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.376412 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 105.730000 0.700000 106.110000 ;
    END
  END EE4END[0]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.5955 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.8236 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 105.59 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 557.143 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 145.990000 0.700000 146.370000 ;
    END
  END E6END[11]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5336 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.7099 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 128.8 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 93.8331 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 490.872 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 144.770000 0.700000 145.150000 ;
    END
  END E6END[10]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.625 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.4032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 85.869 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 458.564 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 143.550000 0.700000 143.930000 ;
    END
  END E6END[9]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.3688 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 93.104 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 48.1831 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 241.527 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.550615 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 141.720000 0.700000 142.100000 ;
    END
  END E6END[8]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.314 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.4938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 213.456 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 156.276 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 815.215 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.85635 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 140.500000 0.700000 140.880000 ;
    END
  END E6END[7]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.32 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 172.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.3258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 30.7463 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 164.109 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 138.670000 0.700000 139.050000 ;
    END
  END E6END[6]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.2356 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.0676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.968 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 103.134 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 522.96 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 137.450000 0.700000 137.830000 ;
    END
  END E6END[5]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.1696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 76.512 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 48.8935 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 243.622 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 135.620000 0.700000 136.000000 ;
    END
  END E6END[4]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.3116 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 124.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1864 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 39.4116 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 207.704 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 134.400000 0.700000 134.780000 ;
    END
  END E6END[3]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.2156 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.2732 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 264.672 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 107.003 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 550.632 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 132.570000 0.700000 132.950000 ;
    END
  END E6END[2]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2174 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.288 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 35.3573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 182.878 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.986768 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 52.7493 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 285.088 LAYER met4  ;
    ANTENNAGATEAREA 1.9125 LAYER met4  ;
    ANTENNAMAXAREACAR 77.5068 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 404.473 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.986768 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 131.350000 0.700000 131.730000 ;
    END
  END E6END[1]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1052 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.16 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met3  ;
    ANTENNAMAXAREACAR 31.0431 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 152.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.691002 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.1838 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 54.784 LAYER met4  ;
    ANTENNAGATEAREA 1.9125 LAYER met4  ;
    ANTENNAMAXAREACAR 36.3679 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 181.149 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.919245 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 130.130000 0.700000 130.510000 ;
    END
  END E6END[0]
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.28 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.174 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 88.820000 0.000000 89.200000 0.700000 ;
    END
  END S1BEG[3]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.145 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 87.440000 0.000000 87.820000 0.700000 ;
    END
  END S1BEG[2]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.871 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 86.060000 0.000000 86.440000 0.700000 ;
    END
  END S1BEG[1]
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.6234 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.009 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 84.220000 0.000000 84.600000 0.700000 ;
    END
  END S1BEG[0]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0218 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.001 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 113.200000 0.000000 113.580000 0.700000 ;
    END
  END S2BEG[7]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.921 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 111.820000 0.000000 112.200000 0.700000 ;
    END
  END S2BEG[6]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.9526 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.537 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 110.440000 0.000000 110.820000 0.700000 ;
    END
  END S2BEG[5]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.599 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 108.600000 0.000000 108.980000 0.700000 ;
    END
  END S2BEG[4]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2982 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.265 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 107.220000 0.000000 107.600000 0.700000 ;
    END
  END S2BEG[3]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1349 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3305 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 105.840000 0.000000 106.220000 0.700000 ;
    END
  END S2BEG[2]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.012 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 104.000000 0.000000 104.380000 0.700000 ;
    END
  END S2BEG[1]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.067 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.227 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 102.620000 0.000000 103.000000 0.700000 ;
    END
  END S2BEG[0]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0602 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.075 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 101.240000 0.000000 101.620000 0.700000 ;
    END
  END S2BEGb[7]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5777 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7805 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.400000 0.000000 99.780000 0.700000 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4578 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.063 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 98.020000 0.000000 98.400000 0.700000 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.07 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 96.640000 0.000000 97.020000 0.700000 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7339 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.4435 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 95.260000 0.000000 95.640000 0.700000 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.0614 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.081 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 93.420000 0.000000 93.800000 0.700000 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.145 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 92.040000 0.000000 92.420000 0.700000 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4006 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.895 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 90.660000 0.000000 91.040000 0.700000 ;
    END
  END S2BEGb[0]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7895 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.7865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.9138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 53.344 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 138.040000 0.000000 138.420000 0.700000 ;
    END
  END S4BEG[15]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7609 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.2098 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 92.256 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 136.200000 0.000000 136.580000 0.700000 ;
    END
  END S4BEG[14]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7814 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.799 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 134.820000 0.000000 135.200000 0.700000 ;
    END
  END S4BEG[13]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4236 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 133.440000 0.000000 133.820000 0.700000 ;
    END
  END S4BEG[12]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0186 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.985 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 131.600000 0.000000 131.980000 0.700000 ;
    END
  END S4BEG[11]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9692 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.62 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 130.220000 0.000000 130.600000 0.700000 ;
    END
  END S4BEG[10]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.599 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 128.840000 0.000000 129.220000 0.700000 ;
    END
  END S4BEG[9]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4482 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.133 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 127.000000 0.000000 127.380000 0.700000 ;
    END
  END S4BEG[8]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.741 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 125.620000 0.000000 126.000000 0.700000 ;
    END
  END S4BEG[7]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0522 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.153 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 124.240000 0.000000 124.620000 0.700000 ;
    END
  END S4BEG[6]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.585 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 122.400000 0.000000 122.780000 0.700000 ;
    END
  END S4BEG[5]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.4621 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.2025 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 121.020000 0.000000 121.400000 0.700000 ;
    END
  END S4BEG[4]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3054 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.419 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 119.640000 0.000000 120.020000 0.700000 ;
    END
  END S4BEG[3]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.741 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 117.800000 0.000000 118.180000 0.700000 ;
    END
  END S4BEG[2]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1288 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.418 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 116.420000 0.000000 116.800000 0.700000 ;
    END
  END S4BEG[1]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.907 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 115.040000 0.000000 115.420000 0.700000 ;
    END
  END S4BEG[0]
  PIN SS4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3786 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.667 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 162.420000 0.000000 162.800000 0.700000 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5568 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.558 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 160.580000 0.000000 160.960000 0.700000 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.051 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 159.200000 0.000000 159.580000 0.700000 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7609 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.5458 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.048 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 157.820000 0.000000 158.200000 0.700000 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 155.980000 0.000000 156.360000 0.700000 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.791 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.729 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 154.600000 0.000000 154.980000 0.700000 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7537 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 153.220000 0.000000 153.600000 0.700000 ;
    END
  END SS4BEG[9]
  PIN SS4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1242 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.395 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 151.380000 0.000000 151.760000 0.700000 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.077 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.159 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.000000 0.000000 150.380000 0.700000 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0419 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.5008 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.808 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 148.620000 0.000000 149.000000 0.700000 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1246 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.397 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 146.780000 0.000000 147.160000 0.700000 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.823 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 145.400000 0.000000 145.780000 0.700000 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3458 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.503 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 144.020000 0.000000 144.400000 0.700000 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.0325 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 142.640000 0.000000 143.020000 0.700000 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.502 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 140.800000 0.000000 141.180000 0.700000 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0218 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.001 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 139.420000 0.000000 139.800000 0.700000 ;
    END
  END SS4BEG[0]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8915 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.1785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.2782 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 142.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.326 LAYER met4  ;
    ANTENNAMAXAREACAR 63.1483 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 322.866 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.831027 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 88.820000 199.560000 89.200000 200.260000 ;
    END
  END S1END[3]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.702 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.123 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 29.9101 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 138.827 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.0684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.16 LAYER met3  ;
    ANTENNAGATEAREA 0.318 LAYER met3  ;
    ANTENNAMAXAREACAR 52.1377 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 258.827 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.700629 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.5876 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 121.408 LAYER met4  ;
    ANTENNAGATEAREA 1.38 LAYER met4  ;
    ANTENNAMAXAREACAR 68.5056 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 346.804 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.942357 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 87.440000 199.560000 87.820000 200.260000 ;
    END
  END S1END[2]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0704 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.083 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 22.8835 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 110.176 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.574 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.528 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 41.0718 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 209.555 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.9366 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 53.936 LAYER met4  ;
    ANTENNAGATEAREA 1.1505 LAYER met4  ;
    ANTENNAMAXAREACAR 49.7085 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 256.435 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 86.060000 199.560000 86.440000 200.260000 ;
    END
  END S1END[1]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.895 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3555 LAYER met2  ;
    ANTENNAMAXAREACAR 11.6007 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 49.0961 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.35757 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.0268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.28 LAYER met3  ;
    ANTENNAGATEAREA 1.1505 LAYER met3  ;
    ANTENNAMAXAREACAR 38.7109 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 187.599 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.515094 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 84.220000 199.560000 84.600000 200.260000 ;
    END
  END S1END[0]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4665 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.1685 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 87.168 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7335 LAYER met4  ;
    ANTENNAMAXAREACAR 54.0151 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 278.161 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 113.200000 199.560000 113.580000 200.260000 ;
    END
  END S2MID[7]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.3814 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 76.209 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6075 LAYER met2  ;
    ANTENNAMAXAREACAR 41.6185 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 198.507 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.606289 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 111.820000 199.560000 112.200000 200.260000 ;
    END
  END S2MID[6]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.219 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 46.7751 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 229.718 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.411 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.992 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 53.9557 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 270.389 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.4448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 120.176 LAYER met4  ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 80.9164 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 414.745 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 110.440000 199.560000 110.820000 200.260000 ;
    END
  END S2MID[5]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3167 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.068 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.496 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.7388 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 66.2784 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 356.768 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.4123 LAYER met4  ;
    ANTENNAMAXAREACAR 56.7203 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 291.751 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.742558 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 108.600000 199.560000 108.980000 200.260000 ;
    END
  END S2MID[4]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 23.7804 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 128.24 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 58.1442 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 305.134 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07583 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 107.220000 199.560000 107.600000 200.260000 ;
    END
  END S2MID[3]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5027 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.0048 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 112.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met4  ;
    ANTENNAMAXAREACAR 45.5889 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 232.768 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.583562 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 105.840000 199.560000 106.220000 200.260000 ;
    END
  END S2MID[2]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.746 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 53.7504 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 287.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7995 LAYER met4  ;
    ANTENNAMAXAREACAR 81.0718 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 426.744 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 104.000000 199.560000 104.380000 200.260000 ;
    END
  END S2MID[1]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4665 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.7388 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 58.2165 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 313.776 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3793 LAYER met4  ;
    ANTENNAMAXAREACAR 47.1819 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 250.903 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 102.620000 199.560000 103.000000 200.260000 ;
    END
  END S2MID[0]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3997 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.333 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.9985 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 96.928 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 78.2434 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 411.98 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 101.240000 199.560000 101.620000 200.260000 ;
    END
  END S2END[7]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.8841 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.9155 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met2  ;
    ANTENNAMAXAREACAR 19.0598 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 87.5167 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.376412 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.992 LAYER met3  ;
    ANTENNAGATEAREA 1.3887 LAYER met3  ;
    ANTENNAMAXAREACAR 25.8059 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 122.485 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.527673 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 99.400000 199.560000 99.780000 200.260000 ;
    END
  END S2END[6]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.3099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.8085 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met2  ;
    ANTENNAMAXAREACAR 31.8501 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 151.831 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.517922 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 32.3815 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 155.285 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.571064 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.9878 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.072 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 38.1335 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 186.301 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 98.020000 199.560000 98.400000 200.260000 ;
    END
  END S2END[5]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.8187 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.6965 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 19.9087 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 80.5003 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 21.7812 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 91.5608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.1808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 198.768 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 48.555 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 241.846 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.748847 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 96.640000 199.560000 97.020000 200.260000 ;
    END
  END S2END[4]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.0302 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.528 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 14.017 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.2792 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.390645 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.515 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.88 LAYER met3  ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 18.2531 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 86.658 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.458019 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.995 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 172.512 LAYER met4  ;
    ANTENNAGATEAREA 1.7067 LAYER met4  ;
    ANTENNAMAXAREACAR 60.0818 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 310.431 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.09371 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 95.260000 199.560000 95.640000 200.260000 ;
    END
  END S2END[3]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0769 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.9975 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 13.6563 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 49.51 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 14.2429 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 53.6692 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.3424 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 141.904 LAYER met4  ;
    ANTENNAGATEAREA 1.7067 LAYER met4  ;
    ANTENNAMAXAREACAR 64.4059 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 322.381 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.695388 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 93.420000 199.560000 93.800000 200.260000 ;
    END
  END S2END[2]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8935 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.0386 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 118.48 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.239 LAYER met4  ;
    ANTENNAMAXAREACAR 42.603 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 214.846 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 92.040000 199.560000 92.420000 200.260000 ;
    END
  END S2END[1]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.2905 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.6305 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met2  ;
    ANTENNAMAXAREACAR 33.2284 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 157.935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.659431 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.574225 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.52 LAYER met3  ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 33.9913 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 162.612 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.712573 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.7513 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 96.08 LAYER met4  ;
    ANTENNAGATEAREA 1.7067 LAYER met4  ;
    ANTENNAMAXAREACAR 81.489 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 418.44 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.857862 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 90.660000 199.560000 91.040000 200.260000 ;
    END
  END S2END[0]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4455 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.0461 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 183.456 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 69.9519 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 372.641 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 138.040000 199.560000 138.420000 200.260000 ;
    END
  END S4END[15]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.2327 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 87.04 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 47.5269 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 247.041 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 136.200000 199.560000 136.580000 200.260000 ;
    END
  END S4END[14]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2427 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.0525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.3928 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 77.232 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 79.4216 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 422.738 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 134.820000 199.560000 135.200000 200.260000 ;
    END
  END S4END[13]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.4446 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.115 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 54.3939 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 268.975 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 133.440000 199.560000 133.820000 200.260000 ;
    END
  END S4END[12]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2141 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.9095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.54 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.0206 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 198.384 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 93.5804 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 487.609 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.67778 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 131.600000 199.560000 131.980000 200.260000 ;
    END
  END S4END[11]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.233 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.939 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 53.317 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 262.99 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 130.220000 199.560000 130.600000 200.260000 ;
    END
  END S4END[10]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.509 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 54.9756 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 271.539 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 128.840000 199.560000 129.220000 200.260000 ;
    END
  END S4END[9]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.683 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.307 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 51.0997 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 252.16 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 127.000000 199.560000 127.380000 200.260000 ;
    END
  END S4END[8]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.5902 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.843 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 57.9252 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 286.288 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 125.620000 199.560000 126.000000 200.260000 ;
    END
  END S4END[7]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8767 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.2225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 23.855 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 121.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 124.240000 199.560000 124.620000 200.260000 ;
    END
  END S4END[6]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.8212 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 111.512 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 51.1831 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 267.277 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 122.400000 199.560000 122.780000 200.260000 ;
    END
  END S4END[5]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0874 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.329 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.4687 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 363.921 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 121.020000 199.560000 121.400000 200.260000 ;
    END
  END S4END[4]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.3744 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.033 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8787 LAYER met2  ;
    ANTENNAMAXAREACAR 21.6041 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 88.9361 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.453458 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.3507 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93 LAYER met3  ;
    ANTENNAGATEAREA 1.3227 LAYER met3  ;
    ANTENNAMAXAREACAR 34.7218 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 159.247 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.498027 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 119.640000 199.560000 120.020000 200.260000 ;
    END
  END S4END[3]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.7041 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.3566 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 136.176 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3227 LAYER met4  ;
    ANTENNAMAXAREACAR 84.0054 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 427.756 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.729603 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 117.800000 199.560000 118.180000 200.260000 ;
    END
  END S4END[2]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6899 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.1705 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 11.674 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.5986 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 14.0228 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 53.1988 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.5274 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 180.224 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 56.1059 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 287.192 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 116.420000 199.560000 116.800000 200.260000 ;
    END
  END S4END[1]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.1678 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.48 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 15.8767 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 64.242 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.5247 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 325.616 LAYER met4  ;
    ANTENNAGATEAREA 1.3557 LAYER met4  ;
    ANTENNAMAXAREACAR 97.0478 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 511.809 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 115.040000 199.560000 115.420000 200.260000 ;
    END
  END S4END[0]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9583 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.5125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.6108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.728 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 73.0341 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 388.234 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 162.420000 199.560000 162.800000 200.260000 ;
    END
  END SS4END[15]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9844 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.761 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.143 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.4778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 72.352 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 72.7621 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 387.303 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 160.580000 199.560000 160.960000 200.260000 ;
    END
  END SS4END[14]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9166 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.422 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.24205 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.9277 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 96.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 36.4412 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 192.157 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 159.200000 199.560000 159.580000 200.260000 ;
    END
  END SS4END[13]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.7474 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.629 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 51.0997 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 252.16 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 157.820000 199.560000 158.200000 200.260000 ;
    END
  END SS4END[12]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9221 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.4495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.8308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 63.568 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 72.8987 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 387.949 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 155.980000 199.560000 156.360000 200.260000 ;
    END
  END SS4END[11]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2499 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.844 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 144.104 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 53.7316 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 284.958 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 154.600000 199.560000 154.980000 200.260000 ;
    END
  END SS4END[10]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7362 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.52 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.056 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.5405 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 185.152 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 91.6104 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 477.291 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 153.220000 199.560000 153.600000 200.260000 ;
    END
  END SS4END[9]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.369 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.737 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 54.0092 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 267.051 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 151.380000 199.560000 151.760000 200.260000 ;
    END
  END SS4END[8]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3849 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.6117 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.728 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 38.1487 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 196.522 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.000000 199.560000 150.380000 200.260000 ;
    END
  END SS4END[7]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3167 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.3275 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 120.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 41.6744 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 220.804 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 148.620000 199.560000 149.000000 200.260000 ;
    END
  END SS4END[6]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.2103 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.7725 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 14.1896 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 52.4247 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 16.697 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 66.8714 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.9658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 80.288 LAYER met4  ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 40.4071 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 194.07 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 146.780000 199.560000 147.160000 200.260000 ;
    END
  END SS4END[5]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.514 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.301 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 7.5758 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.5342 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 8.6547 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 26.3619 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.8588 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 138.384 LAYER met4  ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 49.6224 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 254.914 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 145.400000 199.560000 145.780000 200.260000 ;
    END
  END SS4END[4]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0723 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.9645 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 25.8969 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 110.597 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 26.5156 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 114.811 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.9831 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 167.12 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 82.3241 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 420.782 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 144.020000 199.560000 144.400000 200.260000 ;
    END
  END SS4END[3]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1985 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.4875 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 16.0468 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 72.948 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.532154 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.5466 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99.856 LAYER met3  ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 47.7935 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 239.949 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 142.640000 199.560000 143.020000 200.260000 ;
    END
  END SS4END[2]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.7562 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.857 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met2  ;
    ANTENNAMAXAREACAR 19.0681 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 88.5706 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 140.800000 199.560000 141.180000 200.260000 ;
    END
  END SS4END[1]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7841 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.2975 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 29.02 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 140.164 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 30.1979 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 148.653 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.0433 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 92.304 LAYER met4  ;
    ANTENNAGATEAREA 0.531 LAYER met4  ;
    ANTENNAMAXAREACAR 62.5032 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 322.805 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 139.420000 199.560000 139.800000 200.260000 ;
    END
  END SS4END[0]
  PIN W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 9.350000 0.700000 9.730000 ;
    END
  END W1BEG[3]
  PIN W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 7.520000 0.700000 7.900000 ;
    END
  END W1BEG[2]
  PIN W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.8664 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.616 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 6.300000 0.700000 6.680000 ;
    END
  END W1BEG[1]
  PIN W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 5.080000 0.700000 5.460000 ;
    END
  END W1BEG[0]
  PIN W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 20.940000 0.700000 21.320000 ;
    END
  END W2BEG[7]
  PIN W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.6784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 19.720000 0.700000 20.100000 ;
    END
  END W2BEG[6]
  PIN W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.7965 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.152 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 17.890000 0.700000 18.270000 ;
    END
  END W2BEG[5]
  PIN W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 16.670000 0.700000 17.050000 ;
    END
  END W2BEG[4]
  PIN W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 15.450000 0.700000 15.830000 ;
    END
  END W2BEG[3]
  PIN W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.3548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.096 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 13.620000 0.700000 14.000000 ;
    END
  END W2BEG[2]
  PIN W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.0944 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.832 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 12.400000 0.700000 12.780000 ;
    END
  END W2BEG[1]
  PIN W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 10.570000 0.700000 10.950000 ;
    END
  END W2BEG[0]
  PIN W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.8786 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 143.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 33.140000 0.700000 33.520000 ;
    END
  END W2BEGb[7]
  PIN W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.9174 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 164.888 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 31.310000 0.700000 31.690000 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 30.090000 0.700000 30.470000 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.5995 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.72 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 28.870000 0.700000 29.250000 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 27.040000 0.700000 27.420000 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 25.820000 0.700000 26.200000 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 23.990000 0.700000 24.370000 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 22.770000 0.700000 23.150000 ;
    END
  END W2BEGb[0]
  PIN WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 56.930000 0.700000 57.310000 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 55.100000 0.700000 55.480000 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 53.880000 0.700000 54.260000 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.6444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.432 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 52.660000 0.700000 53.040000 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 50.830000 0.700000 51.210000 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 49.610000 0.700000 49.990000 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 47.780000 0.700000 48.160000 ;
    END
  END WW4BEG[9]
  PIN WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 46.560000 0.700000 46.940000 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.7484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.32 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 44.730000 0.700000 45.110000 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 43.510000 0.700000 43.890000 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 42.290000 0.700000 42.670000 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 40.460000 0.700000 40.840000 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 39.240000 0.700000 39.620000 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 37.410000 0.700000 37.790000 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 36.190000 0.700000 36.570000 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 34.360000 0.700000 34.740000 ;
    END
  END WW4BEG[0]
  PIN W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.4404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 74.620000 0.700000 75.000000 ;
    END
  END W6BEG[11]
  PIN W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 73.400000 0.700000 73.780000 ;
    END
  END W6BEG[10]
  PIN W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 71.570000 0.700000 71.950000 ;
    END
  END W6BEG[9]
  PIN W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.4444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.032 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 70.350000 0.700000 70.730000 ;
    END
  END W6BEG[8]
  PIN W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 68.520000 0.700000 68.900000 ;
    END
  END W6BEG[7]
  PIN W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 67.300000 0.700000 67.680000 ;
    END
  END W6BEG[6]
  PIN W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 66.080000 0.700000 66.460000 ;
    END
  END W6BEG[5]
  PIN W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 64.250000 0.700000 64.630000 ;
    END
  END W6BEG[4]
  PIN W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 63.030000 0.700000 63.410000 ;
    END
  END W6BEG[3]
  PIN W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.5404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.544 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 61.200000 0.700000 61.580000 ;
    END
  END W6BEG[2]
  PIN W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 59.980000 0.700000 60.360000 ;
    END
  END W6BEG[1]
  PIN W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 58.150000 0.700000 58.530000 ;
    END
  END W6BEG[0]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.91292 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.32 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 50.7655 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 262.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.872265 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 30.3315 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 162.704 LAYER met4  ;
    ANTENNAGATEAREA 1.1505 LAYER met4  ;
    ANTENNAMAXAREACAR 77.1293 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 404.4 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.872265 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 9.350000 200.100000 9.730000 ;
    END
  END W1END[3]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.5404 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 256.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1837 LAYER met4  ;
    ANTENNAMAXAREACAR 96.274 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 509.255 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 7.520000 200.100000 7.900000 ;
    END
  END W1END[2]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5874 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 38.7822 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 192.015 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.986768 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.0476 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 86.528 LAYER met4  ;
    ANTENNAGATEAREA 1.1505 LAYER met4  ;
    ANTENNAMAXAREACAR 52.7306 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 267.224 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.986768 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 6.300000 200.100000 6.680000 ;
    END
  END W1END[1]
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 41.2592 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 220.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 59.2053 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 317.168 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1505 LAYER met4  ;
    ANTENNAMAXAREACAR 71.1916 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 369.59 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 5.080000 200.100000 5.460000 ;
    END
  END W1END[0]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2009 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.144 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 100.667 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 502.202 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.0627 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.7996 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.872 LAYER met4  ;
    ANTENNAGATEAREA 0.663 LAYER met4  ;
    ANTENNAMAXAREACAR 104.889 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 526.142 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.36032 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 20.940000 200.100000 21.320000 ;
    END
  END W2MID[7]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.0044 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 139.152 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 69.343 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 349.073 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.6362 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 234.128 LAYER met4  ;
    ANTENNAGATEAREA 1.5882 LAYER met4  ;
    ANTENNAMAXAREACAR 96.8183 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 496.49 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 19.720000 200.100000 20.100000 ;
    END
  END W2MID[6]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.949 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 117.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.2778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.952 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.762 LAYER met4  ;
    ANTENNAMAXAREACAR 46.6336 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 229.252 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.77789 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 17.890000 200.100000 18.270000 ;
    END
  END W2MID[5]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3406 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.2604 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 34.8 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.603 LAYER met4  ;
    ANTENNAMAXAREACAR 57.8684 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 288.542 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.59745 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 16.670000 200.100000 17.050000 ;
    END
  END W2MID[4]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 40.0172 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 213.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.367 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 78.976 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.762 LAYER met4  ;
    ANTENNAMAXAREACAR 37.4385 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 187.73 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 15.450000 200.100000 15.830000 ;
    END
  END W2MID[3]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1496 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.603 LAYER met4  ;
    ANTENNAMAXAREACAR 48.4334 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 235.562 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.540606 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 13.620000 200.100000 14.000000 ;
    END
  END W2MID[2]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.8428 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.432 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.603 LAYER met3  ;
    ANTENNAMAXAREACAR 29.5738 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 150.057 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.606941 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.9826 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.848 LAYER met4  ;
    ANTENNAGATEAREA 0.729 LAYER met4  ;
    ANTENNAMAXAREACAR 33.6651 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 173.168 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 12.400000 200.100000 12.780000 ;
    END
  END W2MID[1]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 30.0444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 160.232 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.603 LAYER met3  ;
    ANTENNAMAXAREACAR 96.3196 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 485.21 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.652843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 10.570000 200.100000 10.950000 ;
    END
  END W2MID[0]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.9764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.336 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7197 LAYER met3  ;
    ANTENNAMAXAREACAR 51.1199 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 242.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.631516 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.9268 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.08 LAYER met4  ;
    ANTENNAGATEAREA 1.0377 LAYER met4  ;
    ANTENNAMAXAREACAR 59.7224 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 289.029 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.631516 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 33.140000 200.100000 33.520000 ;
    END
  END W2END[7]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7866 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 66.2073 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 354.512 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met4  ;
    ANTENNAMAXAREACAR 115.722 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 613.261 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 31.310000 200.100000 31.690000 ;
    END
  END W2END[6]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.3446 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.496 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.3486 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.8 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met4  ;
    ANTENNAMAXAREACAR 49.6302 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 245.902 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 30.090000 200.100000 30.470000 ;
    END
  END W2END[5]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3036 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.2428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.432 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7067 LAYER met4  ;
    ANTENNAMAXAREACAR 56.4286 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 283.138 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.622965 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 28.870000 200.100000 29.250000 ;
    END
  END W2END[4]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5556 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 63.0855 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 339.744 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7997 LAYER met4  ;
    ANTENNAMAXAREACAR 123.728 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 649.524 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.36032 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 27.040000 200.100000 27.420000 ;
    END
  END W2END[3]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.6026 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 141.872 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 70.8199 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 356.119 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.1496 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 135.072 LAYER met4  ;
    ANTENNAGATEAREA 1.5477 LAYER met4  ;
    ANTENNAMAXAREACAR 87.0695 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 443.392 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.80021 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 25.820000 200.100000 26.200000 ;
    END
  END W2END[2]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 38.3299 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 173.991 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.6828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 84.112 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 49.623 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 234.56 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.548637 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 23.990000 200.100000 24.370000 ;
    END
  END W2END[1]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.7346 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 110.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.4097 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0707 LAYER met4  ;
    ANTENNAMAXAREACAR 46.4683 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 235.43 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.653459 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 22.770000 200.100000 23.150000 ;
    END
  END W2END[0]
  PIN WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.544 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 243.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 29.6706 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 149.73 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 56.930000 200.100000 57.310000 ;
    END
  END WW4END[15]
  PIN WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0286 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.1178 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.784 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 91.7944 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 493.468 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 55.100000 200.100000 55.480000 ;
    END
  END WW4END[14]
  PIN WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.8804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 175.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3694 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 29.2294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 156.151 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 53.880000 200.100000 54.260000 ;
    END
  END WW4END[13]
  PIN WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5796 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.9912 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 55.168 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 36.38 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 182.776 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.729187 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 52.660000 200.100000 53.040000 ;
    END
  END WW4END[12]
  PIN WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 42.463 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 226.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.9488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.864 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 30.2222 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 152.718 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 50.830000 200.100000 51.210000 ;
    END
  END WW4END[11]
  PIN WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4186 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.3312 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.648 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 65.7022 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 351.032 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 49.610000 200.100000 49.990000 ;
    END
  END WW4END[10]
  PIN WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.4566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.76 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.8944 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.848 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 72.0169 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 382.742 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 47.780000 200.100000 48.160000 ;
    END
  END WW4END[9]
  PIN WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4076 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.9956 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.584 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 65.8841 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 343.845 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 46.560000 200.100000 46.940000 ;
    END
  END WW4END[8]
  PIN WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8394 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 101.888 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 94.0776 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 487.41 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.67778 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 44.730000 200.100000 45.110000 ;
    END
  END WW4END[7]
  PIN WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.392 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.9236 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.2 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 131.61 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 695.016 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 43.510000 200.100000 43.890000 ;
    END
  END WW4END[6]
  PIN WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.4276 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 114.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.6524 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 58.224 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 53.9118 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 267.732 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.729187 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 42.290000 200.100000 42.670000 ;
    END
  END WW4END[5]
  PIN WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.1364 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.472 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 45.723 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 238.698 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 40.460000 200.100000 40.840000 ;
    END
  END WW4END[4]
  PIN WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.4356 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.6808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.768 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met4  ;
    ANTENNAMAXAREACAR 63.1014 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 325.08 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.502199 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 39.240000 200.100000 39.620000 ;
    END
  END WW4END[3]
  PIN WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.5384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 36.5602 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 166.893 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.7995 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 103.552 LAYER met4  ;
    ANTENNAGATEAREA 0.7527 LAYER met4  ;
    ANTENNAMAXAREACAR 93.2717 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 491.341 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 37.410000 200.100000 37.790000 ;
    END
  END WW4END[2]
  PIN WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 35.8054 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 191.424 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 103.867 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 528.935 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.0372 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.08 LAYER met4  ;
    ANTENNAGATEAREA 0.7527 LAYER met4  ;
    ANTENNAMAXAREACAR 107.902 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 552.955 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.504088 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 36.190000 200.100000 36.570000 ;
    END
  END WW4END[1]
  PIN WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 27.303 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 146.552 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 62.1995 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 313.31 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.449057 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 34.360000 200.100000 34.740000 ;
    END
  END WW4END[0]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.5784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.3698 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 170.128 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 70.3339 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 362.456 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.550615 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 74.620000 200.100000 75.000000 ;
    END
  END W6END[11]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.184 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.8564 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 203.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 86.2781 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 442.786 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.412172 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 73.400000 200.100000 73.780000 ;
    END
  END W6END[10]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 24.7532 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 109.635 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 71.570000 200.100000 71.950000 ;
    END
  END W6END[9]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8276 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.5133 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 180.144 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 68.2951 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 357.03 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 70.350000 200.100000 70.730000 ;
    END
  END W6END[8]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5796 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 62.0853 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 332.528 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 126.98 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 667.765 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 68.520000 200.100000 68.900000 ;
    END
  END W6END[7]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.263 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.0256 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 139.744 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 70.3607 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 362.006 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.550615 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 67.300000 200.100000 67.680000 ;
    END
  END W6END[6]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.3846 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 135.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 23.4532 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 114.571 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 66.080000 200.100000 66.460000 ;
    END
  END W6END[5]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7736 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.7102 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 64.336 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 42.6332 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 209.924 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.796736 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 64.250000 200.100000 64.630000 ;
    END
  END W6END[4]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5796 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.8932 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 49.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 90.5857 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 485.008 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 63.030000 200.100000 63.410000 ;
    END
  END W6END[3]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.9016 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 148.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 19.8008 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 94.4921 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 61.200000 200.100000 61.580000 ;
    END
  END W6END[2]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0774 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 38.7117 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 208.8 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5945 LAYER met4  ;
    ANTENNAMAXAREACAR 87.0588 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 453.777 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 59.980000 200.100000 60.360000 ;
    END
  END W6END[1]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2647 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.872 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 22.0799 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 112.023 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.1971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 66.928 LAYER met4  ;
    ANTENNAGATEAREA 1.6275 LAYER met4  ;
    ANTENNAMAXAREACAR 40.7127 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 198.935 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 58.150000 200.100000 58.530000 ;
    END
  END W6END[0]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2142 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.855 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.0427 LAYER met2  ;
    ANTENNAMAXAREACAR 4.73033 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 5.88282 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.118242 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 163.800000 0.000000 164.180000 0.700000 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1766 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.775 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 163.800000 199.560000 164.180000 200.260000 ;
    END
  END UserCLKo
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.1737 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met3  ;
    ANTENNAMAXAREACAR 36.8626 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 184.874 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.634234 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.4688 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 120.304 LAYER met4  ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 46.7892 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 238.023 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.634234 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 194.180000 0.700000 194.560000 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.101 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.672 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met3  ;
    ANTENNAMAXAREACAR 24.5968 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 119.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.642954 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 31.5306 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 169.104 LAYER met4  ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 43.6524 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 218.82 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 192.350000 0.700000 192.730000 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1576 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.0721 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 220.928 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.193 LAYER met4  ;
    ANTENNAMAXAREACAR 58.2366 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 297.569 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 191.130000 0.700000 191.510000 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.0692 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 145.288 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met3  ;
    ANTENNAMAXAREACAR 77.2696 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 400.914 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.13564 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 46.1502 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 247.536 LAYER met4  ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 97.6585 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 510.274 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.13564 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 189.300000 0.700000 189.680000 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 121.088 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 56.3445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 289.111 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.779245 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 53.2365 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 287.216 LAYER met4  ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 79.864 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 416.001 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 188.080000 0.700000 188.460000 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.7624 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.528 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 47.6926 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 244.567 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.653459 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 35.4318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 191.312 LAYER met4  ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 63.3462 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 329.087 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 186.250000 0.700000 186.630000 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.8022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 106.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.113 LAYER met3  ;
    ANTENNAMAXAREACAR 42.6309 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 214.573 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.689398 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.7581 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 136.272 LAYER met4  ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 53.5689 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 274.777 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 185.030000 0.700000 185.410000 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.3914 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met3  ;
    ANTENNAMAXAREACAR 62.1092 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 317.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.884067 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 37.7973 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 204.864 LAYER met4  ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 78.8078 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 408.243 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 183.200000 0.700000 183.580000 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3429 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.624 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 31.3013 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 163.173 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 69.3828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 372.384 LAYER met4  ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 69.1736 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 357.778 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.09371 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 181.980000 0.700000 182.360000 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.2394 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 98.192 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 56.2469 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 286.289 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.905031 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 65.0757 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 349.888 LAYER met4  ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 84.9969 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 440.868 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 180.760000 0.700000 181.140000 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.3706 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 56.9652 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 307.088 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 84.7851 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 444.803 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 178.930000 0.700000 179.310000 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6572 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.4202 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 89.456 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 57.1447 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 292.499 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.674423 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 177.710000 0.700000 178.090000 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.505 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.16 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met3  ;
    ANTENNAMAXAREACAR 46.134 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 227.854 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.857862 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.2197 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 76.304 LAYER met4  ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 55.6752 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 276.622 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.992502 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 175.880000 0.700000 176.260000 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.9933 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 176.888 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met3  ;
    ANTENNAMAXAREACAR 90.0432 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 469.693 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.939099 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 30.3885 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 164.88 LAYER met4  ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 103.469 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 542.536 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 174.660000 0.700000 175.040000 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.5263 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.064 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 40.0772 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 202.299 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.700629 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 34.749 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 190.032 LAYER met4  ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 84.0198 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 446.291 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 172.830000 0.700000 173.210000 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6836 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 69.5388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 372.736 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 111.745 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 587.758 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.30548 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 171.610000 0.700000 171.990000 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.149 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 79.1289 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 414.412 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 85.6887 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 462.176 LAYER met4  ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 116.986 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 618.598 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 169.780000 0.700000 170.160000 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.232 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met3  ;
    ANTENNAMAXAREACAR 31.4566 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 153.969 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.842138 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 43.3149 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 233.36 LAYER met4  ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 79.7392 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 420.31 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 168.560000 0.700000 168.940000 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.5945 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.824 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 88.5346 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 461.934 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 35.2551 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 189.904 LAYER met4  ;
    ANTENNAGATEAREA 2.193 LAYER met4  ;
    ANTENNAMAXAREACAR 104.611 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 548.529 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.03804 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 167.340000 0.700000 167.720000 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.8839 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.176 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 66.783 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 351.456 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 55.8132 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 299.552 LAYER met4  ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 91.4409 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 483.796 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 165.510000 0.700000 165.890000 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.3214 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.976 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met3  ;
    ANTENNAMAXAREACAR 48.8463 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 249.091 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.884067 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 49.4247 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 266.416 LAYER met4  ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 70.6819 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 366.792 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 164.290000 0.700000 164.670000 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3856 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 63.5541 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 343.184 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.226 LAYER met4  ;
    ANTENNAMAXAREACAR 90.4791 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 476.587 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.2195 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 162.460000 0.700000 162.840000 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.5611 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 179.92 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.113 LAYER met3  ;
    ANTENNAMAXAREACAR 59.854 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 304.614 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.752291 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 60.1491 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 306.395 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.752291 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 161.240000 0.700000 161.620000 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6056 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.304 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1045 LAYER met3  ;
    ANTENNAMAXAREACAR 46.1976 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 226.614 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.609573 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.8846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.992 LAYER met4  ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 47.0302 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 231.47 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 159.410000 0.700000 159.790000 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0094 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.512 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.954 LAYER met3  ;
    ANTENNAMAXAREACAR 24.1245 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 116.49 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 64.7874 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 348.336 LAYER met4  ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 57.6044 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 300.861 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 158.190000 0.700000 158.570000 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.1836 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.888 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.59 LAYER met3  ;
    ANTENNAMAXAREACAR 48.41 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 239.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.757233 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.9799 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 162.24 LAYER met4  ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 61.6549 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 311.381 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 156.360000 0.700000 156.740000 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met3  ;
    ANTENNAMAXAREACAR 29.8262 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 144.927 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 36.7029 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 198.096 LAYER met4  ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 62.511 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 316.061 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 155.140000 0.700000 155.520000 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met3  ;
    ANTENNAMAXAREACAR 41.8898 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 205.277 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.9009 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 247.152 LAYER met4  ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 62.1686 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 314.467 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 153.920000 0.700000 154.300000 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.5946 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 117.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 62.2014 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 327.794 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.886919 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 152.090000 0.700000 152.470000 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.8326 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.4844 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 89.328 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2635 LAYER met4  ;
    ANTENNAMAXAREACAR 51.3654 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 255.39 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 150.870000 0.700000 151.250000 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 70.1434 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 367.645 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.1438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 62.256 LAYER met4  ;
    ANTENNAGATEAREA 2.067 LAYER met4  ;
    ANTENNAMAXAREACAR 85.4859 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 451.66 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 149.040000 0.700000 149.420000 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9606 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.034 LAYER met4  ;
    ANTENNAMAXAREACAR 47.5596 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 233.44 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.98759 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 147.820000 0.700000 148.200000 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 194.180000 200.100000 194.560000 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 192.350000 200.100000 192.730000 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.9884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 191.130000 200.100000 191.510000 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7574 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.368 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 189.300000 200.100000 189.680000 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 188.080000 200.100000 188.460000 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.1834 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 186.250000 200.100000 186.630000 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 185.030000 200.100000 185.410000 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 183.200000 200.100000 183.580000 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 181.980000 200.100000 182.360000 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 180.760000 200.100000 181.140000 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 178.930000 200.100000 179.310000 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 177.710000 200.100000 178.090000 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 175.880000 200.100000 176.260000 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.8174 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 174.660000 200.100000 175.040000 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.0694 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.032 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 172.830000 200.100000 173.210000 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.6784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 171.610000 200.100000 171.990000 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 169.780000 200.100000 170.160000 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 168.560000 200.100000 168.940000 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.4024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.808 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 167.340000 200.100000 167.720000 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 165.510000 200.100000 165.890000 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 164.290000 200.100000 164.670000 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 162.460000 200.100000 162.840000 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 161.240000 200.100000 161.620000 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 159.410000 200.100000 159.790000 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 158.190000 200.100000 158.570000 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.7544 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.352 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 156.360000 200.100000 156.740000 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.5864 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.264 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 155.140000 200.100000 155.520000 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.1104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.016 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 153.920000 200.100000 154.300000 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.0674 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 152.090000 200.100000 152.470000 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.8164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.016 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 150.870000 200.100000 151.250000 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.608 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 149.040000 200.100000 149.420000 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 147.820000 200.100000 148.200000 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6592 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.188 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 53.6193 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 264.674 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 194.160000 0.000000 194.540000 0.700000 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7182 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.483 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 30.3598 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 148.72 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 192.780000 0.000000 193.160000 0.700000 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2299 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 63.1913 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 316.916 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 191.400000 0.000000 191.780000 0.700000 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.7218 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 84.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 40.0865 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 207.227 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.732074 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 190.020000 0.000000 190.400000 0.700000 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8921 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.5258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 88.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 32.5791 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 159.748 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.208175 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 188.180000 0.000000 188.560000 0.700000 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6096 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.94 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 19.9074 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 95.9262 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 186.800000 0.000000 187.180000 0.700000 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.1728 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 81.392 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 37.6199 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 180.369 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.309463 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 185.420000 0.000000 185.800000 0.700000 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8921 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 47.9682 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 257.712 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.9665 LAYER met4  ;
    ANTENNAMAXAREACAR 36.4037 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 180.17 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07583 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 183.580000 0.000000 183.960000 0.700000 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4651 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 55.6848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 299.808 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.214 LAYER met4  ;
    ANTENNAMAXAREACAR 58.8004 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 287.818 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.905577 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 182.200000 0.000000 182.580000 0.700000 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.5873 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 192.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.088 LAYER met2  ;
    ANTENNAMAXAREACAR 25.4346 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 121.195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.614151 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 5.088 LAYER met3  ;
    ANTENNAMAXAREACAR 25.4847 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 121.551 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.622013 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.7588 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 95.184 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 28.8453 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 139.563 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 180.820000 0.000000 181.200000 0.700000 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2983 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.8585 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 54.4158 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 265.796 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.8298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAGATEAREA 0.5145 LAYER met3  ;
    ANTENNAMAXAREACAR 57.9722 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 286.586 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.652588 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.807 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 187.36 LAYER met4  ;
    ANTENNAGATEAREA 5.7192 LAYER met4  ;
    ANTENNAMAXAREACAR 63.8834 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 319.345 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 178.980000 0.000000 179.360000 0.700000 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4159 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.3631 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 34.8162 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 187.568 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 36.492 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 179.802 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.702016 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 177.600000 0.000000 177.980000 0.700000 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.318 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 43.3467 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 234 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 48.1485 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 247.406 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 176.220000 0.000000 176.600000 0.700000 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1235 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.6746 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.056 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.3286 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 77.36 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 27.2482 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 131.831 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 174.380000 0.000000 174.760000 0.700000 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8277 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.9775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 44.1897 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 238.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.214 LAYER met4  ;
    ANTENNAMAXAREACAR 74.5625 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 383.416 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.36032 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 173.000000 0.000000 173.380000 0.700000 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0419 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 89.5287 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 482.176 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.214 LAYER met4  ;
    ANTENNAMAXAREACAR 47.6859 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 246.713 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.36032 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 171.620000 0.000000 172.000000 0.700000 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.09 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.24255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 71.0052 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 382.448 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.214 LAYER met4  ;
    ANTENNAMAXAREACAR 49.4205 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 247.925 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.716691 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 169.780000 0.000000 170.160000 0.700000 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1807 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 71.2509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 382.352 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 42.1857 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 212.794 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.941719 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 168.400000 0.000000 168.780000 0.700000 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0419 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 58.4244 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 313.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.214 LAYER met4  ;
    ANTENNAMAXAREACAR 62.1934 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 317.008 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 167.020000 0.000000 167.400000 0.700000 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.5374 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.542 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met2  ;
    ANTENNAMAXAREACAR 42.3973 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 203.922 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.774004 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3549 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.136 LAYER met3  ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 44.5276 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 216.715 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.89979 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 51.4782 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 278.304 LAYER met4  ;
    ANTENNAGATEAREA 5.214 LAYER met4  ;
    ANTENNAMAXAREACAR 54.4007 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 270.091 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 165.180000 0.000000 165.560000 0.700000 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.064 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.094 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 194.160000 199.560000 194.540000 200.260000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0926 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.237 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 192.780000 199.560000 193.160000 200.260000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.5074 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.311 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 191.400000 199.560000 191.780000 200.260000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9854 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 190.020000 199.560000 190.400000 200.260000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.645 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 188.180000 199.560000 188.560000 200.260000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8088 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.784 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 186.800000 199.560000 187.180000 200.260000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8478 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.131 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 185.420000 199.560000 185.800000 200.260000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.323 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 183.580000 199.560000 183.960000 200.260000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3054 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.419 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 182.200000 199.560000 182.580000 200.260000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7642 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.713 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 180.820000 199.560000 181.200000 200.260000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.543 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.607 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 178.980000 199.560000 179.360000 200.260000 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2242 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.013 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 177.600000 199.560000 177.980000 200.260000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6218 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.001 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 176.220000 199.560000 176.600000 200.260000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1006 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.395 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 174.380000 199.560000 174.760000 200.260000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.6368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 173.000000 199.560000 173.380000 200.260000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.129 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.537 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 171.620000 199.560000 172.000000 200.260000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0194 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.989 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 169.780000 199.560000 170.160000 200.260000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.323 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 168.400000 199.560000 168.780000 200.260000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.1658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.688 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 167.020000 199.560000 167.400000 200.260000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7266 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.407 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 165.180000 199.560000 165.560000 200.260000 ;
    END
  END FrameStrobe_O[0]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 198.900000 195.020000 200.100000 196.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 195.020000 1.200000 196.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.900000 2.850000 200.100000 4.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 1.200000 4.050000 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.070000 199.060000 197.270000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.070000 0.000000 197.270000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 199.060000 4.030000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 0.000000 4.030000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 200.100000 4.050000 ;
        RECT 0.000000 195.020000 200.100000 196.220000 ;
        RECT 2.830000 10.300000 4.030000 10.780000 ;
        RECT 2.830000 4.860000 4.030000 5.340000 ;
        RECT 7.060000 10.300000 8.260000 10.780000 ;
        RECT 7.060000 4.860000 8.260000 5.340000 ;
        RECT 2.830000 15.740000 4.030000 16.220000 ;
        RECT 7.060000 15.740000 8.260000 16.220000 ;
        RECT 2.830000 21.180000 4.030000 21.660000 ;
        RECT 7.060000 21.180000 8.260000 21.660000 ;
        RECT 2.830000 37.500000 4.030000 37.980000 ;
        RECT 7.060000 37.500000 8.260000 37.980000 ;
        RECT 2.830000 32.060000 4.030000 32.540000 ;
        RECT 2.830000 26.620000 4.030000 27.100000 ;
        RECT 7.060000 32.060000 8.260000 32.540000 ;
        RECT 7.060000 26.620000 8.260000 27.100000 ;
        RECT 2.830000 48.380000 4.030000 48.860000 ;
        RECT 2.830000 42.940000 4.030000 43.420000 ;
        RECT 7.060000 48.380000 8.260000 48.860000 ;
        RECT 7.060000 42.940000 8.260000 43.420000 ;
        RECT 52.060000 21.180000 53.260000 21.660000 ;
        RECT 52.060000 15.740000 53.260000 16.220000 ;
        RECT 52.060000 10.300000 53.260000 10.780000 ;
        RECT 52.060000 4.860000 53.260000 5.340000 ;
        RECT 97.060000 21.180000 98.260000 21.660000 ;
        RECT 97.060000 15.740000 98.260000 16.220000 ;
        RECT 97.060000 10.300000 98.260000 10.780000 ;
        RECT 97.060000 4.860000 98.260000 5.340000 ;
        RECT 52.060000 48.380000 53.260000 48.860000 ;
        RECT 52.060000 42.940000 53.260000 43.420000 ;
        RECT 52.060000 37.500000 53.260000 37.980000 ;
        RECT 52.060000 32.060000 53.260000 32.540000 ;
        RECT 52.060000 26.620000 53.260000 27.100000 ;
        RECT 97.060000 48.380000 98.260000 48.860000 ;
        RECT 97.060000 42.940000 98.260000 43.420000 ;
        RECT 97.060000 37.500000 98.260000 37.980000 ;
        RECT 97.060000 32.060000 98.260000 32.540000 ;
        RECT 97.060000 26.620000 98.260000 27.100000 ;
        RECT 2.830000 53.820000 4.030000 54.300000 ;
        RECT 7.060000 53.820000 8.260000 54.300000 ;
        RECT 2.830000 59.260000 4.030000 59.740000 ;
        RECT 7.060000 59.260000 8.260000 59.740000 ;
        RECT 2.830000 70.140000 4.030000 70.620000 ;
        RECT 2.830000 64.700000 4.030000 65.180000 ;
        RECT 7.060000 70.140000 8.260000 70.620000 ;
        RECT 7.060000 64.700000 8.260000 65.180000 ;
        RECT 2.830000 81.020000 4.030000 81.500000 ;
        RECT 7.060000 81.020000 8.260000 81.500000 ;
        RECT 2.830000 75.580000 4.030000 76.060000 ;
        RECT 7.060000 75.580000 8.260000 76.060000 ;
        RECT 2.830000 86.460000 4.030000 86.940000 ;
        RECT 7.060000 86.460000 8.260000 86.940000 ;
        RECT 2.830000 97.340000 4.030000 97.820000 ;
        RECT 2.830000 91.900000 4.030000 92.380000 ;
        RECT 7.060000 97.340000 8.260000 97.820000 ;
        RECT 7.060000 91.900000 8.260000 92.380000 ;
        RECT 52.060000 70.140000 53.260000 70.620000 ;
        RECT 52.060000 64.700000 53.260000 65.180000 ;
        RECT 52.060000 59.260000 53.260000 59.740000 ;
        RECT 52.060000 53.820000 53.260000 54.300000 ;
        RECT 97.060000 70.140000 98.260000 70.620000 ;
        RECT 97.060000 64.700000 98.260000 65.180000 ;
        RECT 97.060000 59.260000 98.260000 59.740000 ;
        RECT 97.060000 53.820000 98.260000 54.300000 ;
        RECT 52.060000 97.340000 53.260000 97.820000 ;
        RECT 52.060000 91.900000 53.260000 92.380000 ;
        RECT 52.060000 86.460000 53.260000 86.940000 ;
        RECT 52.060000 81.020000 53.260000 81.500000 ;
        RECT 52.060000 75.580000 53.260000 76.060000 ;
        RECT 97.060000 97.340000 98.260000 97.820000 ;
        RECT 97.060000 91.900000 98.260000 92.380000 ;
        RECT 97.060000 86.460000 98.260000 86.940000 ;
        RECT 97.060000 81.020000 98.260000 81.500000 ;
        RECT 97.060000 75.580000 98.260000 76.060000 ;
        RECT 142.060000 21.180000 143.260000 21.660000 ;
        RECT 142.060000 15.740000 143.260000 16.220000 ;
        RECT 142.060000 10.300000 143.260000 10.780000 ;
        RECT 142.060000 4.860000 143.260000 5.340000 ;
        RECT 142.060000 48.380000 143.260000 48.860000 ;
        RECT 142.060000 42.940000 143.260000 43.420000 ;
        RECT 142.060000 37.500000 143.260000 37.980000 ;
        RECT 142.060000 32.060000 143.260000 32.540000 ;
        RECT 142.060000 26.620000 143.260000 27.100000 ;
        RECT 196.070000 10.300000 197.270000 10.780000 ;
        RECT 196.070000 4.860000 197.270000 5.340000 ;
        RECT 187.060000 10.300000 188.260000 10.780000 ;
        RECT 187.060000 4.860000 188.260000 5.340000 ;
        RECT 187.060000 21.180000 188.260000 21.660000 ;
        RECT 187.060000 15.740000 188.260000 16.220000 ;
        RECT 196.070000 21.180000 197.270000 21.660000 ;
        RECT 196.070000 15.740000 197.270000 16.220000 ;
        RECT 196.070000 37.500000 197.270000 37.980000 ;
        RECT 187.060000 37.500000 188.260000 37.980000 ;
        RECT 196.070000 32.060000 197.270000 32.540000 ;
        RECT 196.070000 26.620000 197.270000 27.100000 ;
        RECT 187.060000 32.060000 188.260000 32.540000 ;
        RECT 187.060000 26.620000 188.260000 27.100000 ;
        RECT 196.070000 48.380000 197.270000 48.860000 ;
        RECT 196.070000 42.940000 197.270000 43.420000 ;
        RECT 187.060000 48.380000 188.260000 48.860000 ;
        RECT 187.060000 42.940000 188.260000 43.420000 ;
        RECT 142.060000 70.140000 143.260000 70.620000 ;
        RECT 142.060000 64.700000 143.260000 65.180000 ;
        RECT 142.060000 59.260000 143.260000 59.740000 ;
        RECT 142.060000 53.820000 143.260000 54.300000 ;
        RECT 142.060000 97.340000 143.260000 97.820000 ;
        RECT 142.060000 91.900000 143.260000 92.380000 ;
        RECT 142.060000 86.460000 143.260000 86.940000 ;
        RECT 142.060000 81.020000 143.260000 81.500000 ;
        RECT 142.060000 75.580000 143.260000 76.060000 ;
        RECT 187.060000 59.260000 188.260000 59.740000 ;
        RECT 187.060000 53.820000 188.260000 54.300000 ;
        RECT 196.070000 59.260000 197.270000 59.740000 ;
        RECT 196.070000 53.820000 197.270000 54.300000 ;
        RECT 196.070000 70.140000 197.270000 70.620000 ;
        RECT 196.070000 64.700000 197.270000 65.180000 ;
        RECT 187.060000 70.140000 188.260000 70.620000 ;
        RECT 187.060000 64.700000 188.260000 65.180000 ;
        RECT 187.060000 86.460000 188.260000 86.940000 ;
        RECT 187.060000 81.020000 188.260000 81.500000 ;
        RECT 187.060000 75.580000 188.260000 76.060000 ;
        RECT 196.070000 86.460000 197.270000 86.940000 ;
        RECT 196.070000 81.020000 197.270000 81.500000 ;
        RECT 196.070000 75.580000 197.270000 76.060000 ;
        RECT 196.070000 97.340000 197.270000 97.820000 ;
        RECT 196.070000 91.900000 197.270000 92.380000 ;
        RECT 187.060000 97.340000 188.260000 97.820000 ;
        RECT 187.060000 91.900000 188.260000 92.380000 ;
        RECT 2.830000 108.220000 4.030000 108.700000 ;
        RECT 2.830000 102.780000 4.030000 103.260000 ;
        RECT 7.060000 108.220000 8.260000 108.700000 ;
        RECT 7.060000 102.780000 8.260000 103.260000 ;
        RECT 2.830000 113.660000 4.030000 114.140000 ;
        RECT 7.060000 113.660000 8.260000 114.140000 ;
        RECT 2.830000 124.540000 4.030000 125.020000 ;
        RECT 2.830000 119.100000 4.030000 119.580000 ;
        RECT 7.060000 124.540000 8.260000 125.020000 ;
        RECT 7.060000 119.100000 8.260000 119.580000 ;
        RECT 2.830000 135.420000 4.030000 135.900000 ;
        RECT 2.830000 129.980000 4.030000 130.460000 ;
        RECT 7.060000 135.420000 8.260000 135.900000 ;
        RECT 7.060000 129.980000 8.260000 130.460000 ;
        RECT 2.830000 140.860000 4.030000 141.340000 ;
        RECT 7.060000 140.860000 8.260000 141.340000 ;
        RECT 2.830000 146.300000 4.030000 146.780000 ;
        RECT 7.060000 146.300000 8.260000 146.780000 ;
        RECT 52.060000 124.540000 53.260000 125.020000 ;
        RECT 52.060000 119.100000 53.260000 119.580000 ;
        RECT 52.060000 113.660000 53.260000 114.140000 ;
        RECT 52.060000 108.220000 53.260000 108.700000 ;
        RECT 52.060000 102.780000 53.260000 103.260000 ;
        RECT 97.060000 124.540000 98.260000 125.020000 ;
        RECT 97.060000 119.100000 98.260000 119.580000 ;
        RECT 97.060000 113.660000 98.260000 114.140000 ;
        RECT 97.060000 108.220000 98.260000 108.700000 ;
        RECT 97.060000 102.780000 98.260000 103.260000 ;
        RECT 52.060000 146.300000 53.260000 146.780000 ;
        RECT 52.060000 140.860000 53.260000 141.340000 ;
        RECT 52.060000 135.420000 53.260000 135.900000 ;
        RECT 52.060000 129.980000 53.260000 130.460000 ;
        RECT 97.060000 146.300000 98.260000 146.780000 ;
        RECT 97.060000 140.860000 98.260000 141.340000 ;
        RECT 97.060000 135.420000 98.260000 135.900000 ;
        RECT 97.060000 129.980000 98.260000 130.460000 ;
        RECT 2.830000 162.620000 4.030000 163.100000 ;
        RECT 7.060000 162.620000 8.260000 163.100000 ;
        RECT 2.830000 157.180000 4.030000 157.660000 ;
        RECT 2.830000 151.740000 4.030000 152.220000 ;
        RECT 7.060000 157.180000 8.260000 157.660000 ;
        RECT 7.060000 151.740000 8.260000 152.220000 ;
        RECT 2.830000 173.500000 4.030000 173.980000 ;
        RECT 2.830000 168.060000 4.030000 168.540000 ;
        RECT 7.060000 173.500000 8.260000 173.980000 ;
        RECT 7.060000 168.060000 8.260000 168.540000 ;
        RECT 2.830000 178.940000 4.030000 179.420000 ;
        RECT 7.060000 178.940000 8.260000 179.420000 ;
        RECT 2.830000 184.380000 4.030000 184.860000 ;
        RECT 7.060000 184.380000 8.260000 184.860000 ;
        RECT 2.830000 189.820000 4.030000 190.300000 ;
        RECT 7.060000 189.820000 8.260000 190.300000 ;
        RECT 52.060000 173.500000 53.260000 173.980000 ;
        RECT 52.060000 168.060000 53.260000 168.540000 ;
        RECT 52.060000 162.620000 53.260000 163.100000 ;
        RECT 52.060000 157.180000 53.260000 157.660000 ;
        RECT 52.060000 151.740000 53.260000 152.220000 ;
        RECT 97.060000 173.500000 98.260000 173.980000 ;
        RECT 97.060000 168.060000 98.260000 168.540000 ;
        RECT 97.060000 162.620000 98.260000 163.100000 ;
        RECT 97.060000 157.180000 98.260000 157.660000 ;
        RECT 97.060000 151.740000 98.260000 152.220000 ;
        RECT 52.060000 189.820000 53.260000 190.300000 ;
        RECT 52.060000 184.380000 53.260000 184.860000 ;
        RECT 52.060000 178.940000 53.260000 179.420000 ;
        RECT 97.060000 189.820000 98.260000 190.300000 ;
        RECT 97.060000 184.380000 98.260000 184.860000 ;
        RECT 97.060000 178.940000 98.260000 179.420000 ;
        RECT 142.060000 124.540000 143.260000 125.020000 ;
        RECT 142.060000 119.100000 143.260000 119.580000 ;
        RECT 142.060000 113.660000 143.260000 114.140000 ;
        RECT 142.060000 108.220000 143.260000 108.700000 ;
        RECT 142.060000 102.780000 143.260000 103.260000 ;
        RECT 142.060000 146.300000 143.260000 146.780000 ;
        RECT 142.060000 140.860000 143.260000 141.340000 ;
        RECT 142.060000 135.420000 143.260000 135.900000 ;
        RECT 142.060000 129.980000 143.260000 130.460000 ;
        RECT 196.070000 108.220000 197.270000 108.700000 ;
        RECT 196.070000 102.780000 197.270000 103.260000 ;
        RECT 187.060000 108.220000 188.260000 108.700000 ;
        RECT 187.060000 102.780000 188.260000 103.260000 ;
        RECT 187.060000 124.540000 188.260000 125.020000 ;
        RECT 187.060000 119.100000 188.260000 119.580000 ;
        RECT 187.060000 113.660000 188.260000 114.140000 ;
        RECT 196.070000 124.540000 197.270000 125.020000 ;
        RECT 196.070000 119.100000 197.270000 119.580000 ;
        RECT 196.070000 113.660000 197.270000 114.140000 ;
        RECT 196.070000 135.420000 197.270000 135.900000 ;
        RECT 196.070000 129.980000 197.270000 130.460000 ;
        RECT 187.060000 135.420000 188.260000 135.900000 ;
        RECT 187.060000 129.980000 188.260000 130.460000 ;
        RECT 187.060000 146.300000 188.260000 146.780000 ;
        RECT 187.060000 140.860000 188.260000 141.340000 ;
        RECT 196.070000 146.300000 197.270000 146.780000 ;
        RECT 196.070000 140.860000 197.270000 141.340000 ;
        RECT 142.060000 173.500000 143.260000 173.980000 ;
        RECT 142.060000 168.060000 143.260000 168.540000 ;
        RECT 142.060000 162.620000 143.260000 163.100000 ;
        RECT 142.060000 157.180000 143.260000 157.660000 ;
        RECT 142.060000 151.740000 143.260000 152.220000 ;
        RECT 142.060000 189.820000 143.260000 190.300000 ;
        RECT 142.060000 184.380000 143.260000 184.860000 ;
        RECT 142.060000 178.940000 143.260000 179.420000 ;
        RECT 196.070000 162.620000 197.270000 163.100000 ;
        RECT 187.060000 162.620000 188.260000 163.100000 ;
        RECT 196.070000 157.180000 197.270000 157.660000 ;
        RECT 196.070000 151.740000 197.270000 152.220000 ;
        RECT 187.060000 157.180000 188.260000 157.660000 ;
        RECT 187.060000 151.740000 188.260000 152.220000 ;
        RECT 196.070000 173.500000 197.270000 173.980000 ;
        RECT 196.070000 168.060000 197.270000 168.540000 ;
        RECT 187.060000 173.500000 188.260000 173.980000 ;
        RECT 187.060000 168.060000 188.260000 168.540000 ;
        RECT 187.060000 184.380000 188.260000 184.860000 ;
        RECT 187.060000 178.940000 188.260000 179.420000 ;
        RECT 196.070000 184.380000 197.270000 184.860000 ;
        RECT 196.070000 178.940000 197.270000 179.420000 ;
        RECT 196.070000 189.820000 197.270000 190.300000 ;
        RECT 187.060000 189.820000 188.260000 190.300000 ;
      LAYER met4 ;
        RECT 97.060000 2.850000 98.260000 196.220000 ;
        RECT 52.060000 2.850000 53.260000 196.220000 ;
        RECT 7.060000 2.850000 8.260000 196.220000 ;
        RECT 2.830000 0.000000 4.030000 200.260000 ;
        RECT 187.060000 2.850000 188.260000 196.220000 ;
        RECT 142.060000 2.850000 143.260000 196.220000 ;
        RECT 196.070000 0.000000 197.270000 200.260000 ;
    END
# end of P/G power stripe data as pin

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 198.900000 196.820000 200.100000 198.020000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 196.820000 1.200000 198.020000 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.900000 1.050000 200.100000 2.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 1.200000 2.250000 ;
    END
    PORT
      LAYER met4 ;
        RECT 197.870000 199.060000 199.070000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 197.870000 0.000000 199.070000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 199.060000 2.230000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 0.000000 2.230000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 200.100000 2.250000 ;
        RECT 0.000000 196.820000 200.100000 198.020000 ;
        RECT 4.895000 100.060000 6.260000 100.540000 ;
        RECT 50.060000 100.060000 51.260000 100.540000 ;
        RECT 95.060000 100.060000 96.260000 100.540000 ;
        RECT 1.030000 100.060000 2.230000 100.540000 ;
        RECT 140.060000 100.060000 141.260000 100.540000 ;
        RECT 185.060000 100.060000 186.260000 100.540000 ;
        RECT 197.870000 100.060000 199.070000 100.540000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 1.030000 7.580000 2.230000 8.060000 ;
        RECT 1.030000 18.460000 2.230000 18.940000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 1.030000 13.020000 2.230000 13.500000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
        RECT 1.030000 23.900000 2.230000 24.380000 ;
        RECT 4.895000 34.780000 6.260000 35.260000 ;
        RECT 4.895000 29.340000 6.260000 29.820000 ;
        RECT 1.030000 34.780000 2.230000 35.260000 ;
        RECT 1.030000 29.340000 2.230000 29.820000 ;
        RECT 4.895000 45.660000 6.260000 46.140000 ;
        RECT 4.895000 40.220000 6.260000 40.700000 ;
        RECT 1.030000 45.660000 2.230000 46.140000 ;
        RECT 1.030000 40.220000 2.230000 40.700000 ;
        RECT 50.060000 7.580000 51.260000 8.060000 ;
        RECT 50.060000 13.020000 51.260000 13.500000 ;
        RECT 50.060000 18.460000 51.260000 18.940000 ;
        RECT 50.060000 23.900000 51.260000 24.380000 ;
        RECT 95.060000 7.580000 96.260000 8.060000 ;
        RECT 95.060000 13.020000 96.260000 13.500000 ;
        RECT 95.060000 18.460000 96.260000 18.940000 ;
        RECT 95.060000 23.900000 96.260000 24.380000 ;
        RECT 50.060000 29.340000 51.260000 29.820000 ;
        RECT 50.060000 34.780000 51.260000 35.260000 ;
        RECT 50.060000 40.220000 51.260000 40.700000 ;
        RECT 50.060000 45.660000 51.260000 46.140000 ;
        RECT 95.060000 29.340000 96.260000 29.820000 ;
        RECT 95.060000 34.780000 96.260000 35.260000 ;
        RECT 95.060000 40.220000 96.260000 40.700000 ;
        RECT 95.060000 45.660000 96.260000 46.140000 ;
        RECT 1.030000 51.100000 2.230000 51.580000 ;
        RECT 4.895000 51.100000 6.260000 51.580000 ;
        RECT 4.895000 61.980000 6.260000 62.460000 ;
        RECT 4.895000 56.540000 6.260000 57.020000 ;
        RECT 1.030000 56.540000 2.230000 57.020000 ;
        RECT 1.030000 61.980000 2.230000 62.460000 ;
        RECT 4.895000 72.860000 6.260000 73.340000 ;
        RECT 4.895000 67.420000 6.260000 67.900000 ;
        RECT 1.030000 72.860000 2.230000 73.340000 ;
        RECT 1.030000 67.420000 2.230000 67.900000 ;
        RECT 4.895000 78.300000 6.260000 78.780000 ;
        RECT 1.030000 78.300000 2.230000 78.780000 ;
        RECT 4.895000 83.740000 6.260000 84.220000 ;
        RECT 1.030000 83.740000 2.230000 84.220000 ;
        RECT 4.895000 94.620000 6.260000 95.100000 ;
        RECT 4.895000 89.180000 6.260000 89.660000 ;
        RECT 1.030000 94.620000 2.230000 95.100000 ;
        RECT 1.030000 89.180000 2.230000 89.660000 ;
        RECT 50.060000 51.100000 51.260000 51.580000 ;
        RECT 50.060000 56.540000 51.260000 57.020000 ;
        RECT 50.060000 61.980000 51.260000 62.460000 ;
        RECT 50.060000 67.420000 51.260000 67.900000 ;
        RECT 50.060000 72.860000 51.260000 73.340000 ;
        RECT 95.060000 51.100000 96.260000 51.580000 ;
        RECT 95.060000 56.540000 96.260000 57.020000 ;
        RECT 95.060000 61.980000 96.260000 62.460000 ;
        RECT 95.060000 67.420000 96.260000 67.900000 ;
        RECT 95.060000 72.860000 96.260000 73.340000 ;
        RECT 50.060000 78.300000 51.260000 78.780000 ;
        RECT 50.060000 83.740000 51.260000 84.220000 ;
        RECT 50.060000 89.180000 51.260000 89.660000 ;
        RECT 50.060000 94.620000 51.260000 95.100000 ;
        RECT 95.060000 78.300000 96.260000 78.780000 ;
        RECT 95.060000 83.740000 96.260000 84.220000 ;
        RECT 95.060000 89.180000 96.260000 89.660000 ;
        RECT 95.060000 94.620000 96.260000 95.100000 ;
        RECT 140.060000 7.580000 141.260000 8.060000 ;
        RECT 140.060000 13.020000 141.260000 13.500000 ;
        RECT 140.060000 18.460000 141.260000 18.940000 ;
        RECT 140.060000 23.900000 141.260000 24.380000 ;
        RECT 140.060000 29.340000 141.260000 29.820000 ;
        RECT 140.060000 34.780000 141.260000 35.260000 ;
        RECT 140.060000 40.220000 141.260000 40.700000 ;
        RECT 140.060000 45.660000 141.260000 46.140000 ;
        RECT 197.870000 7.580000 199.070000 8.060000 ;
        RECT 185.060000 7.580000 186.260000 8.060000 ;
        RECT 185.060000 23.900000 186.260000 24.380000 ;
        RECT 185.060000 18.460000 186.260000 18.940000 ;
        RECT 185.060000 13.020000 186.260000 13.500000 ;
        RECT 197.870000 13.020000 199.070000 13.500000 ;
        RECT 197.870000 18.460000 199.070000 18.940000 ;
        RECT 197.870000 23.900000 199.070000 24.380000 ;
        RECT 197.870000 34.780000 199.070000 35.260000 ;
        RECT 197.870000 29.340000 199.070000 29.820000 ;
        RECT 185.060000 34.780000 186.260000 35.260000 ;
        RECT 185.060000 29.340000 186.260000 29.820000 ;
        RECT 197.870000 45.660000 199.070000 46.140000 ;
        RECT 197.870000 40.220000 199.070000 40.700000 ;
        RECT 185.060000 45.660000 186.260000 46.140000 ;
        RECT 185.060000 40.220000 186.260000 40.700000 ;
        RECT 140.060000 51.100000 141.260000 51.580000 ;
        RECT 140.060000 56.540000 141.260000 57.020000 ;
        RECT 140.060000 61.980000 141.260000 62.460000 ;
        RECT 140.060000 67.420000 141.260000 67.900000 ;
        RECT 140.060000 72.860000 141.260000 73.340000 ;
        RECT 140.060000 78.300000 141.260000 78.780000 ;
        RECT 140.060000 83.740000 141.260000 84.220000 ;
        RECT 140.060000 89.180000 141.260000 89.660000 ;
        RECT 140.060000 94.620000 141.260000 95.100000 ;
        RECT 185.060000 61.980000 186.260000 62.460000 ;
        RECT 185.060000 56.540000 186.260000 57.020000 ;
        RECT 185.060000 51.100000 186.260000 51.580000 ;
        RECT 197.870000 51.100000 199.070000 51.580000 ;
        RECT 197.870000 56.540000 199.070000 57.020000 ;
        RECT 197.870000 61.980000 199.070000 62.460000 ;
        RECT 197.870000 72.860000 199.070000 73.340000 ;
        RECT 197.870000 67.420000 199.070000 67.900000 ;
        RECT 185.060000 72.860000 186.260000 73.340000 ;
        RECT 185.060000 67.420000 186.260000 67.900000 ;
        RECT 185.060000 78.300000 186.260000 78.780000 ;
        RECT 185.060000 83.740000 186.260000 84.220000 ;
        RECT 197.870000 78.300000 199.070000 78.780000 ;
        RECT 197.870000 83.740000 199.070000 84.220000 ;
        RECT 197.870000 94.620000 199.070000 95.100000 ;
        RECT 197.870000 89.180000 199.070000 89.660000 ;
        RECT 185.060000 94.620000 186.260000 95.100000 ;
        RECT 185.060000 89.180000 186.260000 89.660000 ;
        RECT 4.895000 110.940000 6.260000 111.420000 ;
        RECT 4.895000 105.500000 6.260000 105.980000 ;
        RECT 1.030000 105.500000 2.230000 105.980000 ;
        RECT 1.030000 110.940000 2.230000 111.420000 ;
        RECT 4.895000 116.380000 6.260000 116.860000 ;
        RECT 1.030000 116.380000 2.230000 116.860000 ;
        RECT 4.895000 121.820000 6.260000 122.300000 ;
        RECT 1.030000 121.820000 2.230000 122.300000 ;
        RECT 4.895000 132.700000 6.260000 133.180000 ;
        RECT 1.030000 132.700000 2.230000 133.180000 ;
        RECT 1.030000 127.260000 2.230000 127.740000 ;
        RECT 4.895000 127.260000 6.260000 127.740000 ;
        RECT 1.030000 143.580000 2.230000 144.060000 ;
        RECT 4.895000 143.580000 6.260000 144.060000 ;
        RECT 4.895000 138.140000 6.260000 138.620000 ;
        RECT 1.030000 138.140000 2.230000 138.620000 ;
        RECT 4.895000 149.020000 6.260000 149.500000 ;
        RECT 1.030000 149.020000 2.230000 149.500000 ;
        RECT 50.060000 105.500000 51.260000 105.980000 ;
        RECT 50.060000 110.940000 51.260000 111.420000 ;
        RECT 50.060000 116.380000 51.260000 116.860000 ;
        RECT 50.060000 121.820000 51.260000 122.300000 ;
        RECT 95.060000 105.500000 96.260000 105.980000 ;
        RECT 95.060000 110.940000 96.260000 111.420000 ;
        RECT 95.060000 116.380000 96.260000 116.860000 ;
        RECT 95.060000 121.820000 96.260000 122.300000 ;
        RECT 50.060000 127.260000 51.260000 127.740000 ;
        RECT 50.060000 132.700000 51.260000 133.180000 ;
        RECT 50.060000 138.140000 51.260000 138.620000 ;
        RECT 50.060000 143.580000 51.260000 144.060000 ;
        RECT 50.060000 149.020000 51.260000 149.500000 ;
        RECT 95.060000 127.260000 96.260000 127.740000 ;
        RECT 95.060000 132.700000 96.260000 133.180000 ;
        RECT 95.060000 138.140000 96.260000 138.620000 ;
        RECT 95.060000 143.580000 96.260000 144.060000 ;
        RECT 95.060000 149.020000 96.260000 149.500000 ;
        RECT 4.895000 159.900000 6.260000 160.380000 ;
        RECT 4.895000 154.460000 6.260000 154.940000 ;
        RECT 1.030000 154.460000 2.230000 154.940000 ;
        RECT 1.030000 159.900000 2.230000 160.380000 ;
        RECT 4.895000 170.780000 6.260000 171.260000 ;
        RECT 4.895000 165.340000 6.260000 165.820000 ;
        RECT 1.030000 165.340000 2.230000 165.820000 ;
        RECT 1.030000 170.780000 2.230000 171.260000 ;
        RECT 4.895000 176.220000 6.260000 176.700000 ;
        RECT 1.030000 176.220000 2.230000 176.700000 ;
        RECT 4.895000 187.100000 6.260000 187.580000 ;
        RECT 4.895000 181.660000 6.260000 182.140000 ;
        RECT 1.030000 187.100000 2.230000 187.580000 ;
        RECT 1.030000 181.660000 2.230000 182.140000 ;
        RECT 4.895000 192.540000 6.260000 193.020000 ;
        RECT 1.030000 192.540000 2.230000 193.020000 ;
        RECT 50.060000 154.460000 51.260000 154.940000 ;
        RECT 50.060000 159.900000 51.260000 160.380000 ;
        RECT 50.060000 165.340000 51.260000 165.820000 ;
        RECT 50.060000 170.780000 51.260000 171.260000 ;
        RECT 95.060000 154.460000 96.260000 154.940000 ;
        RECT 95.060000 159.900000 96.260000 160.380000 ;
        RECT 95.060000 165.340000 96.260000 165.820000 ;
        RECT 95.060000 170.780000 96.260000 171.260000 ;
        RECT 50.060000 176.220000 51.260000 176.700000 ;
        RECT 50.060000 181.660000 51.260000 182.140000 ;
        RECT 50.060000 187.100000 51.260000 187.580000 ;
        RECT 50.060000 192.540000 51.260000 193.020000 ;
        RECT 95.060000 176.220000 96.260000 176.700000 ;
        RECT 95.060000 181.660000 96.260000 182.140000 ;
        RECT 95.060000 187.100000 96.260000 187.580000 ;
        RECT 95.060000 192.540000 96.260000 193.020000 ;
        RECT 140.060000 105.500000 141.260000 105.980000 ;
        RECT 140.060000 110.940000 141.260000 111.420000 ;
        RECT 140.060000 116.380000 141.260000 116.860000 ;
        RECT 140.060000 121.820000 141.260000 122.300000 ;
        RECT 140.060000 127.260000 141.260000 127.740000 ;
        RECT 140.060000 132.700000 141.260000 133.180000 ;
        RECT 140.060000 138.140000 141.260000 138.620000 ;
        RECT 140.060000 143.580000 141.260000 144.060000 ;
        RECT 140.060000 149.020000 141.260000 149.500000 ;
        RECT 197.870000 110.940000 199.070000 111.420000 ;
        RECT 197.870000 105.500000 199.070000 105.980000 ;
        RECT 185.060000 105.500000 186.260000 105.980000 ;
        RECT 185.060000 110.940000 186.260000 111.420000 ;
        RECT 185.060000 116.380000 186.260000 116.860000 ;
        RECT 185.060000 121.820000 186.260000 122.300000 ;
        RECT 197.870000 116.380000 199.070000 116.860000 ;
        RECT 197.870000 121.820000 199.070000 122.300000 ;
        RECT 197.870000 132.700000 199.070000 133.180000 ;
        RECT 185.060000 132.700000 186.260000 133.180000 ;
        RECT 185.060000 127.260000 186.260000 127.740000 ;
        RECT 197.870000 127.260000 199.070000 127.740000 ;
        RECT 185.060000 138.140000 186.260000 138.620000 ;
        RECT 185.060000 143.580000 186.260000 144.060000 ;
        RECT 185.060000 149.020000 186.260000 149.500000 ;
        RECT 197.870000 138.140000 199.070000 138.620000 ;
        RECT 197.870000 143.580000 199.070000 144.060000 ;
        RECT 197.870000 149.020000 199.070000 149.500000 ;
        RECT 140.060000 154.460000 141.260000 154.940000 ;
        RECT 140.060000 159.900000 141.260000 160.380000 ;
        RECT 140.060000 165.340000 141.260000 165.820000 ;
        RECT 140.060000 170.780000 141.260000 171.260000 ;
        RECT 140.060000 176.220000 141.260000 176.700000 ;
        RECT 140.060000 181.660000 141.260000 182.140000 ;
        RECT 140.060000 187.100000 141.260000 187.580000 ;
        RECT 140.060000 192.540000 141.260000 193.020000 ;
        RECT 197.870000 159.900000 199.070000 160.380000 ;
        RECT 197.870000 154.460000 199.070000 154.940000 ;
        RECT 185.060000 154.460000 186.260000 154.940000 ;
        RECT 185.060000 159.900000 186.260000 160.380000 ;
        RECT 197.870000 170.780000 199.070000 171.260000 ;
        RECT 197.870000 165.340000 199.070000 165.820000 ;
        RECT 185.060000 165.340000 186.260000 165.820000 ;
        RECT 185.060000 170.780000 186.260000 171.260000 ;
        RECT 185.060000 176.220000 186.260000 176.700000 ;
        RECT 185.060000 181.660000 186.260000 182.140000 ;
        RECT 185.060000 187.100000 186.260000 187.580000 ;
        RECT 197.870000 176.220000 199.070000 176.700000 ;
        RECT 197.870000 181.660000 199.070000 182.140000 ;
        RECT 197.870000 187.100000 199.070000 187.580000 ;
        RECT 197.870000 192.540000 199.070000 193.020000 ;
        RECT 185.060000 192.540000 186.260000 193.020000 ;
      LAYER met4 ;
        RECT 1.030000 0.000000 2.230000 200.260000 ;
        RECT 5.060000 1.050000 6.260000 198.020000 ;
        RECT 50.060000 1.050000 51.260000 198.020000 ;
        RECT 95.060000 1.050000 96.260000 198.020000 ;
        RECT 197.870000 0.000000 199.070000 200.260000 ;
        RECT 140.060000 1.050000 141.260000 198.020000 ;
        RECT 185.060000 1.050000 186.260000 198.020000 ;
        RECT 4.895000 100.060000 6.260000 100.540000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
        RECT 4.895000 34.780000 6.260000 35.260000 ;
        RECT 4.895000 29.340000 6.260000 29.820000 ;
        RECT 4.895000 45.660000 6.260000 46.140000 ;
        RECT 4.895000 40.220000 6.260000 40.700000 ;
        RECT 4.895000 51.100000 6.260000 51.580000 ;
        RECT 4.895000 61.980000 6.260000 62.460000 ;
        RECT 4.895000 56.540000 6.260000 57.020000 ;
        RECT 4.895000 72.860000 6.260000 73.340000 ;
        RECT 4.895000 67.420000 6.260000 67.900000 ;
        RECT 4.895000 78.300000 6.260000 78.780000 ;
        RECT 4.895000 83.740000 6.260000 84.220000 ;
        RECT 4.895000 94.620000 6.260000 95.100000 ;
        RECT 4.895000 89.180000 6.260000 89.660000 ;
        RECT 4.895000 110.940000 6.260000 111.420000 ;
        RECT 4.895000 105.500000 6.260000 105.980000 ;
        RECT 4.895000 116.380000 6.260000 116.860000 ;
        RECT 4.895000 121.820000 6.260000 122.300000 ;
        RECT 4.895000 132.700000 6.260000 133.180000 ;
        RECT 4.895000 127.260000 6.260000 127.740000 ;
        RECT 4.895000 143.580000 6.260000 144.060000 ;
        RECT 4.895000 138.140000 6.260000 138.620000 ;
        RECT 4.895000 149.020000 6.260000 149.500000 ;
        RECT 4.895000 159.900000 6.260000 160.380000 ;
        RECT 4.895000 154.460000 6.260000 154.940000 ;
        RECT 4.895000 170.780000 6.260000 171.260000 ;
        RECT 4.895000 165.340000 6.260000 165.820000 ;
        RECT 4.895000 176.220000 6.260000 176.700000 ;
        RECT 4.895000 187.100000 6.260000 187.580000 ;
        RECT 4.895000 181.660000 6.260000 182.140000 ;
        RECT 4.895000 192.540000 6.260000 193.020000 ;
    END
# end of P/G power stripe data as pin

  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 200.100000 200.260000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 200.100000 200.260000 ;
    LAYER met2 ;
      RECT 194.680000 199.420000 200.100000 200.260000 ;
      RECT 193.300000 199.420000 194.020000 200.260000 ;
      RECT 191.920000 199.420000 192.640000 200.260000 ;
      RECT 190.540000 199.420000 191.260000 200.260000 ;
      RECT 188.700000 199.420000 189.880000 200.260000 ;
      RECT 187.320000 199.420000 188.040000 200.260000 ;
      RECT 185.940000 199.420000 186.660000 200.260000 ;
      RECT 184.100000 199.420000 185.280000 200.260000 ;
      RECT 182.720000 199.420000 183.440000 200.260000 ;
      RECT 181.340000 199.420000 182.060000 200.260000 ;
      RECT 179.500000 199.420000 180.680000 200.260000 ;
      RECT 178.120000 199.420000 178.840000 200.260000 ;
      RECT 176.740000 199.420000 177.460000 200.260000 ;
      RECT 174.900000 199.420000 176.080000 200.260000 ;
      RECT 173.520000 199.420000 174.240000 200.260000 ;
      RECT 172.140000 199.420000 172.860000 200.260000 ;
      RECT 170.300000 199.420000 171.480000 200.260000 ;
      RECT 168.920000 199.420000 169.640000 200.260000 ;
      RECT 167.540000 199.420000 168.260000 200.260000 ;
      RECT 165.700000 199.420000 166.880000 200.260000 ;
      RECT 164.320000 199.420000 165.040000 200.260000 ;
      RECT 162.940000 199.420000 163.660000 200.260000 ;
      RECT 161.100000 199.420000 162.280000 200.260000 ;
      RECT 159.720000 199.420000 160.440000 200.260000 ;
      RECT 158.340000 199.420000 159.060000 200.260000 ;
      RECT 156.500000 199.420000 157.680000 200.260000 ;
      RECT 155.120000 199.420000 155.840000 200.260000 ;
      RECT 153.740000 199.420000 154.460000 200.260000 ;
      RECT 151.900000 199.420000 153.080000 200.260000 ;
      RECT 150.520000 199.420000 151.240000 200.260000 ;
      RECT 149.140000 199.420000 149.860000 200.260000 ;
      RECT 147.300000 199.420000 148.480000 200.260000 ;
      RECT 145.920000 199.420000 146.640000 200.260000 ;
      RECT 144.540000 199.420000 145.260000 200.260000 ;
      RECT 143.160000 199.420000 143.880000 200.260000 ;
      RECT 141.320000 199.420000 142.500000 200.260000 ;
      RECT 139.940000 199.420000 140.660000 200.260000 ;
      RECT 138.560000 199.420000 139.280000 200.260000 ;
      RECT 136.720000 199.420000 137.900000 200.260000 ;
      RECT 135.340000 199.420000 136.060000 200.260000 ;
      RECT 133.960000 199.420000 134.680000 200.260000 ;
      RECT 132.120000 199.420000 133.300000 200.260000 ;
      RECT 130.740000 199.420000 131.460000 200.260000 ;
      RECT 129.360000 199.420000 130.080000 200.260000 ;
      RECT 127.520000 199.420000 128.700000 200.260000 ;
      RECT 126.140000 199.420000 126.860000 200.260000 ;
      RECT 124.760000 199.420000 125.480000 200.260000 ;
      RECT 122.920000 199.420000 124.100000 200.260000 ;
      RECT 121.540000 199.420000 122.260000 200.260000 ;
      RECT 120.160000 199.420000 120.880000 200.260000 ;
      RECT 118.320000 199.420000 119.500000 200.260000 ;
      RECT 116.940000 199.420000 117.660000 200.260000 ;
      RECT 115.560000 199.420000 116.280000 200.260000 ;
      RECT 113.720000 199.420000 114.900000 200.260000 ;
      RECT 112.340000 199.420000 113.060000 200.260000 ;
      RECT 110.960000 199.420000 111.680000 200.260000 ;
      RECT 109.120000 199.420000 110.300000 200.260000 ;
      RECT 107.740000 199.420000 108.460000 200.260000 ;
      RECT 106.360000 199.420000 107.080000 200.260000 ;
      RECT 104.520000 199.420000 105.700000 200.260000 ;
      RECT 103.140000 199.420000 103.860000 200.260000 ;
      RECT 101.760000 199.420000 102.480000 200.260000 ;
      RECT 99.920000 199.420000 101.100000 200.260000 ;
      RECT 98.540000 199.420000 99.260000 200.260000 ;
      RECT 97.160000 199.420000 97.880000 200.260000 ;
      RECT 95.780000 199.420000 96.500000 200.260000 ;
      RECT 93.940000 199.420000 95.120000 200.260000 ;
      RECT 92.560000 199.420000 93.280000 200.260000 ;
      RECT 91.180000 199.420000 91.900000 200.260000 ;
      RECT 89.340000 199.420000 90.520000 200.260000 ;
      RECT 87.960000 199.420000 88.680000 200.260000 ;
      RECT 86.580000 199.420000 87.300000 200.260000 ;
      RECT 84.740000 199.420000 85.920000 200.260000 ;
      RECT 83.360000 199.420000 84.080000 200.260000 ;
      RECT 81.980000 199.420000 82.700000 200.260000 ;
      RECT 80.140000 199.420000 81.320000 200.260000 ;
      RECT 78.760000 199.420000 79.480000 200.260000 ;
      RECT 77.380000 199.420000 78.100000 200.260000 ;
      RECT 75.540000 199.420000 76.720000 200.260000 ;
      RECT 74.160000 199.420000 74.880000 200.260000 ;
      RECT 72.780000 199.420000 73.500000 200.260000 ;
      RECT 70.940000 199.420000 72.120000 200.260000 ;
      RECT 69.560000 199.420000 70.280000 200.260000 ;
      RECT 68.180000 199.420000 68.900000 200.260000 ;
      RECT 66.340000 199.420000 67.520000 200.260000 ;
      RECT 64.960000 199.420000 65.680000 200.260000 ;
      RECT 63.580000 199.420000 64.300000 200.260000 ;
      RECT 61.740000 199.420000 62.920000 200.260000 ;
      RECT 60.360000 199.420000 61.080000 200.260000 ;
      RECT 58.980000 199.420000 59.700000 200.260000 ;
      RECT 57.140000 199.420000 58.320000 200.260000 ;
      RECT 55.760000 199.420000 56.480000 200.260000 ;
      RECT 54.380000 199.420000 55.100000 200.260000 ;
      RECT 53.000000 199.420000 53.720000 200.260000 ;
      RECT 51.160000 199.420000 52.340000 200.260000 ;
      RECT 49.780000 199.420000 50.500000 200.260000 ;
      RECT 48.400000 199.420000 49.120000 200.260000 ;
      RECT 46.560000 199.420000 47.740000 200.260000 ;
      RECT 45.180000 199.420000 45.900000 200.260000 ;
      RECT 43.800000 199.420000 44.520000 200.260000 ;
      RECT 41.960000 199.420000 43.140000 200.260000 ;
      RECT 40.580000 199.420000 41.300000 200.260000 ;
      RECT 39.200000 199.420000 39.920000 200.260000 ;
      RECT 37.360000 199.420000 38.540000 200.260000 ;
      RECT 35.980000 199.420000 36.700000 200.260000 ;
      RECT 34.600000 199.420000 35.320000 200.260000 ;
      RECT 32.760000 199.420000 33.940000 200.260000 ;
      RECT 31.380000 199.420000 32.100000 200.260000 ;
      RECT 30.000000 199.420000 30.720000 200.260000 ;
      RECT 28.160000 199.420000 29.340000 200.260000 ;
      RECT 26.780000 199.420000 27.500000 200.260000 ;
      RECT 25.400000 199.420000 26.120000 200.260000 ;
      RECT 23.560000 199.420000 24.740000 200.260000 ;
      RECT 22.180000 199.420000 22.900000 200.260000 ;
      RECT 20.800000 199.420000 21.520000 200.260000 ;
      RECT 18.960000 199.420000 20.140000 200.260000 ;
      RECT 17.580000 199.420000 18.300000 200.260000 ;
      RECT 16.200000 199.420000 16.920000 200.260000 ;
      RECT 14.360000 199.420000 15.540000 200.260000 ;
      RECT 12.980000 199.420000 13.700000 200.260000 ;
      RECT 11.600000 199.420000 12.320000 200.260000 ;
      RECT 9.760000 199.420000 10.940000 200.260000 ;
      RECT 8.380000 199.420000 9.100000 200.260000 ;
      RECT 7.000000 199.420000 7.720000 200.260000 ;
      RECT 5.620000 199.420000 6.340000 200.260000 ;
      RECT 0.000000 199.420000 4.960000 200.260000 ;
      RECT 0.000000 0.840000 200.100000 199.420000 ;
      RECT 194.680000 0.000000 200.100000 0.840000 ;
      RECT 193.300000 0.000000 194.020000 0.840000 ;
      RECT 191.920000 0.000000 192.640000 0.840000 ;
      RECT 190.540000 0.000000 191.260000 0.840000 ;
      RECT 188.700000 0.000000 189.880000 0.840000 ;
      RECT 187.320000 0.000000 188.040000 0.840000 ;
      RECT 185.940000 0.000000 186.660000 0.840000 ;
      RECT 184.100000 0.000000 185.280000 0.840000 ;
      RECT 182.720000 0.000000 183.440000 0.840000 ;
      RECT 181.340000 0.000000 182.060000 0.840000 ;
      RECT 179.500000 0.000000 180.680000 0.840000 ;
      RECT 178.120000 0.000000 178.840000 0.840000 ;
      RECT 176.740000 0.000000 177.460000 0.840000 ;
      RECT 174.900000 0.000000 176.080000 0.840000 ;
      RECT 173.520000 0.000000 174.240000 0.840000 ;
      RECT 172.140000 0.000000 172.860000 0.840000 ;
      RECT 170.300000 0.000000 171.480000 0.840000 ;
      RECT 168.920000 0.000000 169.640000 0.840000 ;
      RECT 167.540000 0.000000 168.260000 0.840000 ;
      RECT 165.700000 0.000000 166.880000 0.840000 ;
      RECT 164.320000 0.000000 165.040000 0.840000 ;
      RECT 162.940000 0.000000 163.660000 0.840000 ;
      RECT 161.100000 0.000000 162.280000 0.840000 ;
      RECT 159.720000 0.000000 160.440000 0.840000 ;
      RECT 158.340000 0.000000 159.060000 0.840000 ;
      RECT 156.500000 0.000000 157.680000 0.840000 ;
      RECT 155.120000 0.000000 155.840000 0.840000 ;
      RECT 153.740000 0.000000 154.460000 0.840000 ;
      RECT 151.900000 0.000000 153.080000 0.840000 ;
      RECT 150.520000 0.000000 151.240000 0.840000 ;
      RECT 149.140000 0.000000 149.860000 0.840000 ;
      RECT 147.300000 0.000000 148.480000 0.840000 ;
      RECT 145.920000 0.000000 146.640000 0.840000 ;
      RECT 144.540000 0.000000 145.260000 0.840000 ;
      RECT 143.160000 0.000000 143.880000 0.840000 ;
      RECT 141.320000 0.000000 142.500000 0.840000 ;
      RECT 139.940000 0.000000 140.660000 0.840000 ;
      RECT 138.560000 0.000000 139.280000 0.840000 ;
      RECT 136.720000 0.000000 137.900000 0.840000 ;
      RECT 135.340000 0.000000 136.060000 0.840000 ;
      RECT 133.960000 0.000000 134.680000 0.840000 ;
      RECT 132.120000 0.000000 133.300000 0.840000 ;
      RECT 130.740000 0.000000 131.460000 0.840000 ;
      RECT 129.360000 0.000000 130.080000 0.840000 ;
      RECT 127.520000 0.000000 128.700000 0.840000 ;
      RECT 126.140000 0.000000 126.860000 0.840000 ;
      RECT 124.760000 0.000000 125.480000 0.840000 ;
      RECT 122.920000 0.000000 124.100000 0.840000 ;
      RECT 121.540000 0.000000 122.260000 0.840000 ;
      RECT 120.160000 0.000000 120.880000 0.840000 ;
      RECT 118.320000 0.000000 119.500000 0.840000 ;
      RECT 116.940000 0.000000 117.660000 0.840000 ;
      RECT 115.560000 0.000000 116.280000 0.840000 ;
      RECT 113.720000 0.000000 114.900000 0.840000 ;
      RECT 112.340000 0.000000 113.060000 0.840000 ;
      RECT 110.960000 0.000000 111.680000 0.840000 ;
      RECT 109.120000 0.000000 110.300000 0.840000 ;
      RECT 107.740000 0.000000 108.460000 0.840000 ;
      RECT 106.360000 0.000000 107.080000 0.840000 ;
      RECT 104.520000 0.000000 105.700000 0.840000 ;
      RECT 103.140000 0.000000 103.860000 0.840000 ;
      RECT 101.760000 0.000000 102.480000 0.840000 ;
      RECT 99.920000 0.000000 101.100000 0.840000 ;
      RECT 98.540000 0.000000 99.260000 0.840000 ;
      RECT 97.160000 0.000000 97.880000 0.840000 ;
      RECT 95.780000 0.000000 96.500000 0.840000 ;
      RECT 93.940000 0.000000 95.120000 0.840000 ;
      RECT 92.560000 0.000000 93.280000 0.840000 ;
      RECT 91.180000 0.000000 91.900000 0.840000 ;
      RECT 89.340000 0.000000 90.520000 0.840000 ;
      RECT 87.960000 0.000000 88.680000 0.840000 ;
      RECT 86.580000 0.000000 87.300000 0.840000 ;
      RECT 84.740000 0.000000 85.920000 0.840000 ;
      RECT 83.360000 0.000000 84.080000 0.840000 ;
      RECT 81.980000 0.000000 82.700000 0.840000 ;
      RECT 80.140000 0.000000 81.320000 0.840000 ;
      RECT 78.760000 0.000000 79.480000 0.840000 ;
      RECT 77.380000 0.000000 78.100000 0.840000 ;
      RECT 75.540000 0.000000 76.720000 0.840000 ;
      RECT 74.160000 0.000000 74.880000 0.840000 ;
      RECT 72.780000 0.000000 73.500000 0.840000 ;
      RECT 70.940000 0.000000 72.120000 0.840000 ;
      RECT 69.560000 0.000000 70.280000 0.840000 ;
      RECT 68.180000 0.000000 68.900000 0.840000 ;
      RECT 66.340000 0.000000 67.520000 0.840000 ;
      RECT 64.960000 0.000000 65.680000 0.840000 ;
      RECT 63.580000 0.000000 64.300000 0.840000 ;
      RECT 61.740000 0.000000 62.920000 0.840000 ;
      RECT 60.360000 0.000000 61.080000 0.840000 ;
      RECT 58.980000 0.000000 59.700000 0.840000 ;
      RECT 57.140000 0.000000 58.320000 0.840000 ;
      RECT 55.760000 0.000000 56.480000 0.840000 ;
      RECT 54.380000 0.000000 55.100000 0.840000 ;
      RECT 53.000000 0.000000 53.720000 0.840000 ;
      RECT 51.160000 0.000000 52.340000 0.840000 ;
      RECT 49.780000 0.000000 50.500000 0.840000 ;
      RECT 48.400000 0.000000 49.120000 0.840000 ;
      RECT 46.560000 0.000000 47.740000 0.840000 ;
      RECT 45.180000 0.000000 45.900000 0.840000 ;
      RECT 43.800000 0.000000 44.520000 0.840000 ;
      RECT 41.960000 0.000000 43.140000 0.840000 ;
      RECT 40.580000 0.000000 41.300000 0.840000 ;
      RECT 39.200000 0.000000 39.920000 0.840000 ;
      RECT 37.360000 0.000000 38.540000 0.840000 ;
      RECT 35.980000 0.000000 36.700000 0.840000 ;
      RECT 34.600000 0.000000 35.320000 0.840000 ;
      RECT 32.760000 0.000000 33.940000 0.840000 ;
      RECT 31.380000 0.000000 32.100000 0.840000 ;
      RECT 30.000000 0.000000 30.720000 0.840000 ;
      RECT 28.160000 0.000000 29.340000 0.840000 ;
      RECT 26.780000 0.000000 27.500000 0.840000 ;
      RECT 25.400000 0.000000 26.120000 0.840000 ;
      RECT 23.560000 0.000000 24.740000 0.840000 ;
      RECT 22.180000 0.000000 22.900000 0.840000 ;
      RECT 20.800000 0.000000 21.520000 0.840000 ;
      RECT 18.960000 0.000000 20.140000 0.840000 ;
      RECT 17.580000 0.000000 18.300000 0.840000 ;
      RECT 16.200000 0.000000 16.920000 0.840000 ;
      RECT 14.360000 0.000000 15.540000 0.840000 ;
      RECT 12.980000 0.000000 13.700000 0.840000 ;
      RECT 11.600000 0.000000 12.320000 0.840000 ;
      RECT 9.760000 0.000000 10.940000 0.840000 ;
      RECT 8.380000 0.000000 9.100000 0.840000 ;
      RECT 7.000000 0.000000 7.720000 0.840000 ;
      RECT 5.620000 0.000000 6.340000 0.840000 ;
      RECT 0.000000 0.000000 4.960000 0.840000 ;
    LAYER met3 ;
      RECT 0.000000 198.320000 200.100000 200.260000 ;
      RECT 1.000000 193.880000 199.100000 194.720000 ;
      RECT 0.000000 193.320000 200.100000 193.880000 ;
      RECT 199.370000 193.030000 200.100000 193.320000 ;
      RECT 0.000000 193.030000 0.730000 193.320000 ;
      RECT 186.560000 192.240000 197.570000 193.320000 ;
      RECT 141.560000 192.240000 184.760000 193.320000 ;
      RECT 96.560000 192.240000 139.760000 193.320000 ;
      RECT 51.560000 192.240000 94.760000 193.320000 ;
      RECT 6.560000 192.240000 49.760000 193.320000 ;
      RECT 2.530000 192.240000 4.595000 193.320000 ;
      RECT 1.000000 192.050000 199.100000 192.240000 ;
      RECT 0.000000 191.810000 200.100000 192.050000 ;
      RECT 1.000000 190.830000 199.100000 191.810000 ;
      RECT 0.000000 190.600000 200.100000 190.830000 ;
      RECT 197.570000 189.980000 200.100000 190.600000 ;
      RECT 0.000000 189.980000 2.530000 190.600000 ;
      RECT 197.570000 189.520000 199.100000 189.980000 ;
      RECT 188.560000 189.520000 195.770000 190.600000 ;
      RECT 143.560000 189.520000 186.760000 190.600000 ;
      RECT 98.560000 189.520000 141.760000 190.600000 ;
      RECT 53.560000 189.520000 96.760000 190.600000 ;
      RECT 8.560000 189.520000 51.760000 190.600000 ;
      RECT 4.330000 189.520000 6.760000 190.600000 ;
      RECT 1.000000 189.520000 2.530000 189.980000 ;
      RECT 1.000000 189.000000 199.100000 189.520000 ;
      RECT 0.000000 188.760000 200.100000 189.000000 ;
      RECT 1.000000 187.880000 199.100000 188.760000 ;
      RECT 199.370000 186.930000 200.100000 187.780000 ;
      RECT 0.000000 186.930000 0.730000 187.780000 ;
      RECT 186.560000 186.800000 197.570000 187.880000 ;
      RECT 141.560000 186.800000 184.760000 187.880000 ;
      RECT 96.560000 186.800000 139.760000 187.880000 ;
      RECT 51.560000 186.800000 94.760000 187.880000 ;
      RECT 6.560000 186.800000 49.760000 187.880000 ;
      RECT 2.530000 186.800000 4.595000 187.880000 ;
      RECT 1.000000 185.950000 199.100000 186.800000 ;
      RECT 0.000000 185.710000 200.100000 185.950000 ;
      RECT 1.000000 185.160000 199.100000 185.710000 ;
      RECT 197.570000 184.730000 199.100000 185.160000 ;
      RECT 1.000000 184.730000 2.530000 185.160000 ;
      RECT 197.570000 184.080000 200.100000 184.730000 ;
      RECT 188.560000 184.080000 195.770000 185.160000 ;
      RECT 143.560000 184.080000 186.760000 185.160000 ;
      RECT 98.560000 184.080000 141.760000 185.160000 ;
      RECT 53.560000 184.080000 96.760000 185.160000 ;
      RECT 8.560000 184.080000 51.760000 185.160000 ;
      RECT 4.330000 184.080000 6.760000 185.160000 ;
      RECT 0.000000 184.080000 2.530000 184.730000 ;
      RECT 0.000000 183.880000 200.100000 184.080000 ;
      RECT 1.000000 182.900000 199.100000 183.880000 ;
      RECT 0.000000 182.660000 200.100000 182.900000 ;
      RECT 1.000000 182.440000 199.100000 182.660000 ;
      RECT 199.370000 181.440000 200.100000 181.680000 ;
      RECT 0.000000 181.440000 0.730000 181.680000 ;
      RECT 186.560000 181.360000 197.570000 182.440000 ;
      RECT 141.560000 181.360000 184.760000 182.440000 ;
      RECT 96.560000 181.360000 139.760000 182.440000 ;
      RECT 51.560000 181.360000 94.760000 182.440000 ;
      RECT 6.560000 181.360000 49.760000 182.440000 ;
      RECT 2.530000 181.360000 4.595000 182.440000 ;
      RECT 1.000000 180.460000 199.100000 181.360000 ;
      RECT 0.000000 179.720000 200.100000 180.460000 ;
      RECT 197.570000 179.610000 200.100000 179.720000 ;
      RECT 0.000000 179.610000 2.530000 179.720000 ;
      RECT 197.570000 178.640000 199.100000 179.610000 ;
      RECT 188.560000 178.640000 195.770000 179.720000 ;
      RECT 143.560000 178.640000 186.760000 179.720000 ;
      RECT 98.560000 178.640000 141.760000 179.720000 ;
      RECT 53.560000 178.640000 96.760000 179.720000 ;
      RECT 8.560000 178.640000 51.760000 179.720000 ;
      RECT 4.330000 178.640000 6.760000 179.720000 ;
      RECT 1.000000 178.640000 2.530000 179.610000 ;
      RECT 1.000000 178.630000 199.100000 178.640000 ;
      RECT 0.000000 178.390000 200.100000 178.630000 ;
      RECT 1.000000 177.410000 199.100000 178.390000 ;
      RECT 0.000000 177.000000 200.100000 177.410000 ;
      RECT 199.370000 176.560000 200.100000 177.000000 ;
      RECT 0.000000 176.560000 0.730000 177.000000 ;
      RECT 186.560000 175.920000 197.570000 177.000000 ;
      RECT 141.560000 175.920000 184.760000 177.000000 ;
      RECT 96.560000 175.920000 139.760000 177.000000 ;
      RECT 51.560000 175.920000 94.760000 177.000000 ;
      RECT 6.560000 175.920000 49.760000 177.000000 ;
      RECT 2.530000 175.920000 4.595000 177.000000 ;
      RECT 1.000000 175.580000 199.100000 175.920000 ;
      RECT 0.000000 175.340000 200.100000 175.580000 ;
      RECT 1.000000 174.360000 199.100000 175.340000 ;
      RECT 0.000000 174.280000 200.100000 174.360000 ;
      RECT 197.570000 173.510000 200.100000 174.280000 ;
      RECT 0.000000 173.510000 2.530000 174.280000 ;
      RECT 197.570000 173.200000 199.100000 173.510000 ;
      RECT 188.560000 173.200000 195.770000 174.280000 ;
      RECT 143.560000 173.200000 186.760000 174.280000 ;
      RECT 98.560000 173.200000 141.760000 174.280000 ;
      RECT 53.560000 173.200000 96.760000 174.280000 ;
      RECT 8.560000 173.200000 51.760000 174.280000 ;
      RECT 4.330000 173.200000 6.760000 174.280000 ;
      RECT 1.000000 173.200000 2.530000 173.510000 ;
      RECT 1.000000 172.530000 199.100000 173.200000 ;
      RECT 0.000000 172.290000 200.100000 172.530000 ;
      RECT 1.000000 171.560000 199.100000 172.290000 ;
      RECT 199.370000 170.480000 200.100000 171.310000 ;
      RECT 186.560000 170.480000 197.570000 171.560000 ;
      RECT 141.560000 170.480000 184.760000 171.560000 ;
      RECT 96.560000 170.480000 139.760000 171.560000 ;
      RECT 51.560000 170.480000 94.760000 171.560000 ;
      RECT 6.560000 170.480000 49.760000 171.560000 ;
      RECT 2.530000 170.480000 4.595000 171.560000 ;
      RECT 0.000000 170.480000 0.730000 171.310000 ;
      RECT 0.000000 170.460000 200.100000 170.480000 ;
      RECT 1.000000 169.480000 199.100000 170.460000 ;
      RECT 0.000000 169.240000 200.100000 169.480000 ;
      RECT 1.000000 168.840000 199.100000 169.240000 ;
      RECT 197.570000 168.260000 199.100000 168.840000 ;
      RECT 1.000000 168.260000 2.530000 168.840000 ;
      RECT 197.570000 168.020000 200.100000 168.260000 ;
      RECT 0.000000 168.020000 2.530000 168.260000 ;
      RECT 197.570000 167.760000 199.100000 168.020000 ;
      RECT 188.560000 167.760000 195.770000 168.840000 ;
      RECT 143.560000 167.760000 186.760000 168.840000 ;
      RECT 98.560000 167.760000 141.760000 168.840000 ;
      RECT 53.560000 167.760000 96.760000 168.840000 ;
      RECT 8.560000 167.760000 51.760000 168.840000 ;
      RECT 4.330000 167.760000 6.760000 168.840000 ;
      RECT 1.000000 167.760000 2.530000 168.020000 ;
      RECT 1.000000 167.040000 199.100000 167.760000 ;
      RECT 0.000000 166.190000 200.100000 167.040000 ;
      RECT 1.000000 166.120000 199.100000 166.190000 ;
      RECT 199.370000 165.040000 200.100000 165.210000 ;
      RECT 186.560000 165.040000 197.570000 166.120000 ;
      RECT 141.560000 165.040000 184.760000 166.120000 ;
      RECT 96.560000 165.040000 139.760000 166.120000 ;
      RECT 51.560000 165.040000 94.760000 166.120000 ;
      RECT 6.560000 165.040000 49.760000 166.120000 ;
      RECT 2.530000 165.040000 4.595000 166.120000 ;
      RECT 0.000000 165.040000 0.730000 165.210000 ;
      RECT 0.000000 164.970000 200.100000 165.040000 ;
      RECT 1.000000 163.990000 199.100000 164.970000 ;
      RECT 0.000000 163.400000 200.100000 163.990000 ;
      RECT 197.570000 163.140000 200.100000 163.400000 ;
      RECT 0.000000 163.140000 2.530000 163.400000 ;
      RECT 197.570000 162.320000 199.100000 163.140000 ;
      RECT 188.560000 162.320000 195.770000 163.400000 ;
      RECT 143.560000 162.320000 186.760000 163.400000 ;
      RECT 98.560000 162.320000 141.760000 163.400000 ;
      RECT 53.560000 162.320000 96.760000 163.400000 ;
      RECT 8.560000 162.320000 51.760000 163.400000 ;
      RECT 4.330000 162.320000 6.760000 163.400000 ;
      RECT 1.000000 162.320000 2.530000 163.140000 ;
      RECT 1.000000 162.160000 199.100000 162.320000 ;
      RECT 0.000000 161.920000 200.100000 162.160000 ;
      RECT 1.000000 160.940000 199.100000 161.920000 ;
      RECT 0.000000 160.680000 200.100000 160.940000 ;
      RECT 199.370000 160.090000 200.100000 160.680000 ;
      RECT 0.000000 160.090000 0.730000 160.680000 ;
      RECT 186.560000 159.600000 197.570000 160.680000 ;
      RECT 141.560000 159.600000 184.760000 160.680000 ;
      RECT 96.560000 159.600000 139.760000 160.680000 ;
      RECT 51.560000 159.600000 94.760000 160.680000 ;
      RECT 6.560000 159.600000 49.760000 160.680000 ;
      RECT 2.530000 159.600000 4.595000 160.680000 ;
      RECT 1.000000 159.110000 199.100000 159.600000 ;
      RECT 0.000000 158.870000 200.100000 159.110000 ;
      RECT 1.000000 157.960000 199.100000 158.870000 ;
      RECT 197.570000 157.890000 199.100000 157.960000 ;
      RECT 1.000000 157.890000 2.530000 157.960000 ;
      RECT 197.570000 157.040000 200.100000 157.890000 ;
      RECT 0.000000 157.040000 2.530000 157.890000 ;
      RECT 197.570000 156.880000 199.100000 157.040000 ;
      RECT 188.560000 156.880000 195.770000 157.960000 ;
      RECT 143.560000 156.880000 186.760000 157.960000 ;
      RECT 98.560000 156.880000 141.760000 157.960000 ;
      RECT 53.560000 156.880000 96.760000 157.960000 ;
      RECT 8.560000 156.880000 51.760000 157.960000 ;
      RECT 4.330000 156.880000 6.760000 157.960000 ;
      RECT 1.000000 156.880000 2.530000 157.040000 ;
      RECT 1.000000 156.060000 199.100000 156.880000 ;
      RECT 0.000000 155.820000 200.100000 156.060000 ;
      RECT 1.000000 155.240000 199.100000 155.820000 ;
      RECT 199.370000 154.600000 200.100000 154.840000 ;
      RECT 0.000000 154.600000 0.730000 154.840000 ;
      RECT 186.560000 154.160000 197.570000 155.240000 ;
      RECT 141.560000 154.160000 184.760000 155.240000 ;
      RECT 96.560000 154.160000 139.760000 155.240000 ;
      RECT 51.560000 154.160000 94.760000 155.240000 ;
      RECT 6.560000 154.160000 49.760000 155.240000 ;
      RECT 2.530000 154.160000 4.595000 155.240000 ;
      RECT 1.000000 153.620000 199.100000 154.160000 ;
      RECT 0.000000 152.770000 200.100000 153.620000 ;
      RECT 1.000000 152.520000 199.100000 152.770000 ;
      RECT 197.570000 151.790000 199.100000 152.520000 ;
      RECT 1.000000 151.790000 2.530000 152.520000 ;
      RECT 197.570000 151.550000 200.100000 151.790000 ;
      RECT 0.000000 151.550000 2.530000 151.790000 ;
      RECT 197.570000 151.440000 199.100000 151.550000 ;
      RECT 188.560000 151.440000 195.770000 152.520000 ;
      RECT 143.560000 151.440000 186.760000 152.520000 ;
      RECT 98.560000 151.440000 141.760000 152.520000 ;
      RECT 53.560000 151.440000 96.760000 152.520000 ;
      RECT 8.560000 151.440000 51.760000 152.520000 ;
      RECT 4.330000 151.440000 6.760000 152.520000 ;
      RECT 1.000000 151.440000 2.530000 151.550000 ;
      RECT 1.000000 150.570000 199.100000 151.440000 ;
      RECT 0.000000 149.800000 200.100000 150.570000 ;
      RECT 199.370000 149.720000 200.100000 149.800000 ;
      RECT 0.000000 149.720000 0.730000 149.800000 ;
      RECT 199.370000 148.720000 200.100000 148.740000 ;
      RECT 186.560000 148.720000 197.570000 149.800000 ;
      RECT 141.560000 148.720000 184.760000 149.800000 ;
      RECT 96.560000 148.720000 139.760000 149.800000 ;
      RECT 51.560000 148.720000 94.760000 149.800000 ;
      RECT 6.560000 148.720000 49.760000 149.800000 ;
      RECT 2.530000 148.720000 4.595000 149.800000 ;
      RECT 0.000000 148.720000 0.730000 148.740000 ;
      RECT 0.000000 148.500000 200.100000 148.720000 ;
      RECT 1.000000 147.520000 199.100000 148.500000 ;
      RECT 0.000000 147.080000 200.100000 147.520000 ;
      RECT 197.570000 146.670000 200.100000 147.080000 ;
      RECT 0.000000 146.670000 2.530000 147.080000 ;
      RECT 197.570000 146.000000 199.100000 146.670000 ;
      RECT 188.560000 146.000000 195.770000 147.080000 ;
      RECT 143.560000 146.000000 186.760000 147.080000 ;
      RECT 98.560000 146.000000 141.760000 147.080000 ;
      RECT 53.560000 146.000000 96.760000 147.080000 ;
      RECT 8.560000 146.000000 51.760000 147.080000 ;
      RECT 4.330000 146.000000 6.760000 147.080000 ;
      RECT 1.000000 146.000000 2.530000 146.670000 ;
      RECT 1.000000 145.690000 199.100000 146.000000 ;
      RECT 0.000000 145.450000 200.100000 145.690000 ;
      RECT 1.000000 144.470000 199.100000 145.450000 ;
      RECT 0.000000 144.360000 200.100000 144.470000 ;
      RECT 199.370000 144.230000 200.100000 144.360000 ;
      RECT 0.000000 144.230000 0.730000 144.360000 ;
      RECT 186.560000 143.280000 197.570000 144.360000 ;
      RECT 141.560000 143.280000 184.760000 144.360000 ;
      RECT 96.560000 143.280000 139.760000 144.360000 ;
      RECT 51.560000 143.280000 94.760000 144.360000 ;
      RECT 6.560000 143.280000 49.760000 144.360000 ;
      RECT 2.530000 143.280000 4.595000 144.360000 ;
      RECT 1.000000 143.250000 199.100000 143.280000 ;
      RECT 0.000000 142.400000 200.100000 143.250000 ;
      RECT 1.000000 141.640000 199.100000 142.400000 ;
      RECT 197.570000 141.420000 199.100000 141.640000 ;
      RECT 1.000000 141.420000 2.530000 141.640000 ;
      RECT 197.570000 141.180000 200.100000 141.420000 ;
      RECT 0.000000 141.180000 2.530000 141.420000 ;
      RECT 197.570000 140.560000 199.100000 141.180000 ;
      RECT 188.560000 140.560000 195.770000 141.640000 ;
      RECT 143.560000 140.560000 186.760000 141.640000 ;
      RECT 98.560000 140.560000 141.760000 141.640000 ;
      RECT 53.560000 140.560000 96.760000 141.640000 ;
      RECT 8.560000 140.560000 51.760000 141.640000 ;
      RECT 4.330000 140.560000 6.760000 141.640000 ;
      RECT 1.000000 140.560000 2.530000 141.180000 ;
      RECT 1.000000 140.200000 199.100000 140.560000 ;
      RECT 0.000000 139.350000 200.100000 140.200000 ;
      RECT 1.000000 138.920000 199.100000 139.350000 ;
      RECT 199.370000 138.130000 200.100000 138.370000 ;
      RECT 0.000000 138.130000 0.730000 138.370000 ;
      RECT 186.560000 137.840000 197.570000 138.920000 ;
      RECT 141.560000 137.840000 184.760000 138.920000 ;
      RECT 96.560000 137.840000 139.760000 138.920000 ;
      RECT 51.560000 137.840000 94.760000 138.920000 ;
      RECT 6.560000 137.840000 49.760000 138.920000 ;
      RECT 2.530000 137.840000 4.595000 138.920000 ;
      RECT 1.000000 137.150000 199.100000 137.840000 ;
      RECT 0.000000 136.300000 200.100000 137.150000 ;
      RECT 1.000000 136.200000 199.100000 136.300000 ;
      RECT 197.570000 135.320000 199.100000 136.200000 ;
      RECT 1.000000 135.320000 2.530000 136.200000 ;
      RECT 197.570000 135.120000 200.100000 135.320000 ;
      RECT 188.560000 135.120000 195.770000 136.200000 ;
      RECT 143.560000 135.120000 186.760000 136.200000 ;
      RECT 98.560000 135.120000 141.760000 136.200000 ;
      RECT 53.560000 135.120000 96.760000 136.200000 ;
      RECT 8.560000 135.120000 51.760000 136.200000 ;
      RECT 4.330000 135.120000 6.760000 136.200000 ;
      RECT 0.000000 135.120000 2.530000 135.320000 ;
      RECT 0.000000 135.080000 200.100000 135.120000 ;
      RECT 1.000000 134.100000 199.100000 135.080000 ;
      RECT 0.000000 133.480000 200.100000 134.100000 ;
      RECT 199.370000 133.250000 200.100000 133.480000 ;
      RECT 0.000000 133.250000 0.730000 133.480000 ;
      RECT 186.560000 132.400000 197.570000 133.480000 ;
      RECT 141.560000 132.400000 184.760000 133.480000 ;
      RECT 96.560000 132.400000 139.760000 133.480000 ;
      RECT 51.560000 132.400000 94.760000 133.480000 ;
      RECT 6.560000 132.400000 49.760000 133.480000 ;
      RECT 2.530000 132.400000 4.595000 133.480000 ;
      RECT 1.000000 132.270000 199.100000 132.400000 ;
      RECT 0.000000 132.030000 200.100000 132.270000 ;
      RECT 1.000000 131.050000 199.100000 132.030000 ;
      RECT 0.000000 130.810000 200.100000 131.050000 ;
      RECT 1.000000 130.760000 199.100000 130.810000 ;
      RECT 197.570000 129.830000 199.100000 130.760000 ;
      RECT 1.000000 129.830000 2.530000 130.760000 ;
      RECT 197.570000 129.680000 200.100000 129.830000 ;
      RECT 188.560000 129.680000 195.770000 130.760000 ;
      RECT 143.560000 129.680000 186.760000 130.760000 ;
      RECT 98.560000 129.680000 141.760000 130.760000 ;
      RECT 53.560000 129.680000 96.760000 130.760000 ;
      RECT 8.560000 129.680000 51.760000 130.760000 ;
      RECT 4.330000 129.680000 6.760000 130.760000 ;
      RECT 0.000000 129.680000 2.530000 129.830000 ;
      RECT 0.000000 128.980000 200.100000 129.680000 ;
      RECT 1.000000 128.040000 199.100000 128.980000 ;
      RECT 199.370000 127.760000 200.100000 128.000000 ;
      RECT 0.000000 127.760000 0.730000 128.000000 ;
      RECT 186.560000 126.960000 197.570000 128.040000 ;
      RECT 141.560000 126.960000 184.760000 128.040000 ;
      RECT 96.560000 126.960000 139.760000 128.040000 ;
      RECT 51.560000 126.960000 94.760000 128.040000 ;
      RECT 6.560000 126.960000 49.760000 128.040000 ;
      RECT 2.530000 126.960000 4.595000 128.040000 ;
      RECT 1.000000 126.780000 199.100000 126.960000 ;
      RECT 0.000000 125.930000 200.100000 126.780000 ;
      RECT 1.000000 125.320000 199.100000 125.930000 ;
      RECT 197.570000 124.950000 199.100000 125.320000 ;
      RECT 1.000000 124.950000 2.530000 125.320000 ;
      RECT 197.570000 124.710000 200.100000 124.950000 ;
      RECT 0.000000 124.710000 2.530000 124.950000 ;
      RECT 197.570000 124.240000 199.100000 124.710000 ;
      RECT 188.560000 124.240000 195.770000 125.320000 ;
      RECT 143.560000 124.240000 186.760000 125.320000 ;
      RECT 98.560000 124.240000 141.760000 125.320000 ;
      RECT 53.560000 124.240000 96.760000 125.320000 ;
      RECT 8.560000 124.240000 51.760000 125.320000 ;
      RECT 4.330000 124.240000 6.760000 125.320000 ;
      RECT 1.000000 124.240000 2.530000 124.710000 ;
      RECT 1.000000 123.730000 199.100000 124.240000 ;
      RECT 0.000000 122.880000 200.100000 123.730000 ;
      RECT 1.000000 122.600000 199.100000 122.880000 ;
      RECT 199.370000 121.660000 200.100000 121.900000 ;
      RECT 0.000000 121.660000 0.730000 121.900000 ;
      RECT 186.560000 121.520000 197.570000 122.600000 ;
      RECT 141.560000 121.520000 184.760000 122.600000 ;
      RECT 96.560000 121.520000 139.760000 122.600000 ;
      RECT 51.560000 121.520000 94.760000 122.600000 ;
      RECT 6.560000 121.520000 49.760000 122.600000 ;
      RECT 2.530000 121.520000 4.595000 122.600000 ;
      RECT 1.000000 120.680000 199.100000 121.520000 ;
      RECT 0.000000 119.880000 200.100000 120.680000 ;
      RECT 197.570000 119.830000 200.100000 119.880000 ;
      RECT 0.000000 119.830000 2.530000 119.880000 ;
      RECT 197.570000 118.850000 199.100000 119.830000 ;
      RECT 1.000000 118.850000 2.530000 119.830000 ;
      RECT 197.570000 118.800000 200.100000 118.850000 ;
      RECT 188.560000 118.800000 195.770000 119.880000 ;
      RECT 143.560000 118.800000 186.760000 119.880000 ;
      RECT 98.560000 118.800000 141.760000 119.880000 ;
      RECT 53.560000 118.800000 96.760000 119.880000 ;
      RECT 8.560000 118.800000 51.760000 119.880000 ;
      RECT 4.330000 118.800000 6.760000 119.880000 ;
      RECT 0.000000 118.800000 2.530000 118.850000 ;
      RECT 0.000000 118.610000 200.100000 118.800000 ;
      RECT 1.000000 117.630000 199.100000 118.610000 ;
      RECT 0.000000 117.390000 200.100000 117.630000 ;
      RECT 1.000000 117.160000 199.100000 117.390000 ;
      RECT 199.370000 116.080000 200.100000 116.410000 ;
      RECT 186.560000 116.080000 197.570000 117.160000 ;
      RECT 141.560000 116.080000 184.760000 117.160000 ;
      RECT 96.560000 116.080000 139.760000 117.160000 ;
      RECT 51.560000 116.080000 94.760000 117.160000 ;
      RECT 6.560000 116.080000 49.760000 117.160000 ;
      RECT 2.530000 116.080000 4.595000 117.160000 ;
      RECT 0.000000 116.080000 0.730000 116.410000 ;
      RECT 0.000000 115.560000 200.100000 116.080000 ;
      RECT 1.000000 114.580000 199.100000 115.560000 ;
      RECT 0.000000 114.440000 200.100000 114.580000 ;
      RECT 197.570000 114.340000 200.100000 114.440000 ;
      RECT 0.000000 114.340000 2.530000 114.440000 ;
      RECT 197.570000 113.360000 199.100000 114.340000 ;
      RECT 188.560000 113.360000 195.770000 114.440000 ;
      RECT 143.560000 113.360000 186.760000 114.440000 ;
      RECT 98.560000 113.360000 141.760000 114.440000 ;
      RECT 53.560000 113.360000 96.760000 114.440000 ;
      RECT 8.560000 113.360000 51.760000 114.440000 ;
      RECT 4.330000 113.360000 6.760000 114.440000 ;
      RECT 1.000000 113.360000 2.530000 114.340000 ;
      RECT 0.000000 112.510000 200.100000 113.360000 ;
      RECT 1.000000 111.720000 199.100000 112.510000 ;
      RECT 199.370000 111.290000 200.100000 111.530000 ;
      RECT 0.000000 111.290000 0.730000 111.530000 ;
      RECT 186.560000 110.640000 197.570000 111.720000 ;
      RECT 141.560000 110.640000 184.760000 111.720000 ;
      RECT 96.560000 110.640000 139.760000 111.720000 ;
      RECT 51.560000 110.640000 94.760000 111.720000 ;
      RECT 6.560000 110.640000 49.760000 111.720000 ;
      RECT 2.530000 110.640000 4.595000 111.720000 ;
      RECT 1.000000 110.310000 199.100000 110.640000 ;
      RECT 0.000000 109.460000 200.100000 110.310000 ;
      RECT 1.000000 109.000000 199.100000 109.460000 ;
      RECT 197.570000 108.480000 199.100000 109.000000 ;
      RECT 1.000000 108.480000 2.530000 109.000000 ;
      RECT 197.570000 108.240000 200.100000 108.480000 ;
      RECT 0.000000 108.240000 2.530000 108.480000 ;
      RECT 197.570000 107.920000 199.100000 108.240000 ;
      RECT 188.560000 107.920000 195.770000 109.000000 ;
      RECT 143.560000 107.920000 186.760000 109.000000 ;
      RECT 98.560000 107.920000 141.760000 109.000000 ;
      RECT 53.560000 107.920000 96.760000 109.000000 ;
      RECT 8.560000 107.920000 51.760000 109.000000 ;
      RECT 4.330000 107.920000 6.760000 109.000000 ;
      RECT 1.000000 107.920000 2.530000 108.240000 ;
      RECT 1.000000 107.260000 199.100000 107.920000 ;
      RECT 0.000000 106.410000 200.100000 107.260000 ;
      RECT 1.000000 106.280000 199.100000 106.410000 ;
      RECT 199.370000 105.200000 200.100000 105.430000 ;
      RECT 186.560000 105.200000 197.570000 106.280000 ;
      RECT 141.560000 105.200000 184.760000 106.280000 ;
      RECT 96.560000 105.200000 139.760000 106.280000 ;
      RECT 51.560000 105.200000 94.760000 106.280000 ;
      RECT 6.560000 105.200000 49.760000 106.280000 ;
      RECT 2.530000 105.200000 4.595000 106.280000 ;
      RECT 0.000000 105.200000 0.730000 105.430000 ;
      RECT 0.000000 105.190000 200.100000 105.200000 ;
      RECT 1.000000 104.210000 199.100000 105.190000 ;
      RECT 0.000000 103.970000 200.100000 104.210000 ;
      RECT 1.000000 103.560000 199.100000 103.970000 ;
      RECT 197.570000 102.990000 199.100000 103.560000 ;
      RECT 1.000000 102.990000 2.530000 103.560000 ;
      RECT 197.570000 102.480000 200.100000 102.990000 ;
      RECT 188.560000 102.480000 195.770000 103.560000 ;
      RECT 143.560000 102.480000 186.760000 103.560000 ;
      RECT 98.560000 102.480000 141.760000 103.560000 ;
      RECT 53.560000 102.480000 96.760000 103.560000 ;
      RECT 8.560000 102.480000 51.760000 103.560000 ;
      RECT 4.330000 102.480000 6.760000 103.560000 ;
      RECT 0.000000 102.480000 2.530000 102.990000 ;
      RECT 0.000000 102.140000 200.100000 102.480000 ;
      RECT 1.000000 101.160000 199.100000 102.140000 ;
      RECT 0.000000 100.920000 200.100000 101.160000 ;
      RECT 1.000000 100.840000 199.100000 100.920000 ;
      RECT 199.370000 99.760000 200.100000 99.940000 ;
      RECT 186.560000 99.760000 197.570000 100.840000 ;
      RECT 141.560000 99.760000 184.760000 100.840000 ;
      RECT 96.560000 99.760000 139.760000 100.840000 ;
      RECT 51.560000 99.760000 94.760000 100.840000 ;
      RECT 6.560000 99.760000 49.760000 100.840000 ;
      RECT 2.530000 99.760000 4.595000 100.840000 ;
      RECT 0.000000 99.760000 0.730000 99.940000 ;
      RECT 0.000000 99.090000 200.100000 99.760000 ;
      RECT 1.000000 98.120000 199.100000 99.090000 ;
      RECT 197.570000 98.110000 199.100000 98.120000 ;
      RECT 1.000000 98.110000 2.530000 98.120000 ;
      RECT 197.570000 97.870000 200.100000 98.110000 ;
      RECT 0.000000 97.870000 2.530000 98.110000 ;
      RECT 197.570000 97.040000 199.100000 97.870000 ;
      RECT 188.560000 97.040000 195.770000 98.120000 ;
      RECT 143.560000 97.040000 186.760000 98.120000 ;
      RECT 98.560000 97.040000 141.760000 98.120000 ;
      RECT 53.560000 97.040000 96.760000 98.120000 ;
      RECT 8.560000 97.040000 51.760000 98.120000 ;
      RECT 4.330000 97.040000 6.760000 98.120000 ;
      RECT 1.000000 97.040000 2.530000 97.870000 ;
      RECT 1.000000 96.890000 199.100000 97.040000 ;
      RECT 0.000000 96.040000 200.100000 96.890000 ;
      RECT 1.000000 95.400000 199.100000 96.040000 ;
      RECT 199.370000 94.820000 200.100000 95.060000 ;
      RECT 0.000000 94.820000 0.730000 95.060000 ;
      RECT 186.560000 94.320000 197.570000 95.400000 ;
      RECT 141.560000 94.320000 184.760000 95.400000 ;
      RECT 96.560000 94.320000 139.760000 95.400000 ;
      RECT 51.560000 94.320000 94.760000 95.400000 ;
      RECT 6.560000 94.320000 49.760000 95.400000 ;
      RECT 2.530000 94.320000 4.595000 95.400000 ;
      RECT 1.000000 93.840000 199.100000 94.320000 ;
      RECT 0.000000 93.600000 200.100000 93.840000 ;
      RECT 1.000000 92.680000 199.100000 93.600000 ;
      RECT 197.570000 92.620000 199.100000 92.680000 ;
      RECT 1.000000 92.620000 2.530000 92.680000 ;
      RECT 197.570000 91.770000 200.100000 92.620000 ;
      RECT 0.000000 91.770000 2.530000 92.620000 ;
      RECT 197.570000 91.600000 199.100000 91.770000 ;
      RECT 188.560000 91.600000 195.770000 92.680000 ;
      RECT 143.560000 91.600000 186.760000 92.680000 ;
      RECT 98.560000 91.600000 141.760000 92.680000 ;
      RECT 53.560000 91.600000 96.760000 92.680000 ;
      RECT 8.560000 91.600000 51.760000 92.680000 ;
      RECT 4.330000 91.600000 6.760000 92.680000 ;
      RECT 1.000000 91.600000 2.530000 91.770000 ;
      RECT 1.000000 90.790000 199.100000 91.600000 ;
      RECT 0.000000 90.550000 200.100000 90.790000 ;
      RECT 1.000000 89.960000 199.100000 90.550000 ;
      RECT 199.370000 88.880000 200.100000 89.570000 ;
      RECT 186.560000 88.880000 197.570000 89.960000 ;
      RECT 141.560000 88.880000 184.760000 89.960000 ;
      RECT 96.560000 88.880000 139.760000 89.960000 ;
      RECT 51.560000 88.880000 94.760000 89.960000 ;
      RECT 6.560000 88.880000 49.760000 89.960000 ;
      RECT 2.530000 88.880000 4.595000 89.960000 ;
      RECT 0.000000 88.880000 0.730000 89.570000 ;
      RECT 0.000000 88.720000 200.100000 88.880000 ;
      RECT 1.000000 87.740000 199.100000 88.720000 ;
      RECT 0.000000 87.500000 200.100000 87.740000 ;
      RECT 1.000000 87.240000 199.100000 87.500000 ;
      RECT 197.570000 86.520000 199.100000 87.240000 ;
      RECT 1.000000 86.520000 2.530000 87.240000 ;
      RECT 197.570000 86.160000 200.100000 86.520000 ;
      RECT 188.560000 86.160000 195.770000 87.240000 ;
      RECT 143.560000 86.160000 186.760000 87.240000 ;
      RECT 98.560000 86.160000 141.760000 87.240000 ;
      RECT 53.560000 86.160000 96.760000 87.240000 ;
      RECT 8.560000 86.160000 51.760000 87.240000 ;
      RECT 4.330000 86.160000 6.760000 87.240000 ;
      RECT 0.000000 86.160000 2.530000 86.520000 ;
      RECT 0.000000 85.670000 200.100000 86.160000 ;
      RECT 1.000000 84.690000 199.100000 85.670000 ;
      RECT 0.000000 84.520000 200.100000 84.690000 ;
      RECT 199.370000 84.450000 200.100000 84.520000 ;
      RECT 0.000000 84.450000 0.730000 84.520000 ;
      RECT 199.370000 83.440000 200.100000 83.470000 ;
      RECT 186.560000 83.440000 197.570000 84.520000 ;
      RECT 141.560000 83.440000 184.760000 84.520000 ;
      RECT 96.560000 83.440000 139.760000 84.520000 ;
      RECT 51.560000 83.440000 94.760000 84.520000 ;
      RECT 6.560000 83.440000 49.760000 84.520000 ;
      RECT 2.530000 83.440000 4.595000 84.520000 ;
      RECT 0.000000 83.440000 0.730000 83.470000 ;
      RECT 0.000000 82.620000 200.100000 83.440000 ;
      RECT 1.000000 81.800000 199.100000 82.620000 ;
      RECT 197.570000 81.640000 199.100000 81.800000 ;
      RECT 1.000000 81.640000 2.530000 81.800000 ;
      RECT 197.570000 81.400000 200.100000 81.640000 ;
      RECT 0.000000 81.400000 2.530000 81.640000 ;
      RECT 197.570000 80.720000 199.100000 81.400000 ;
      RECT 188.560000 80.720000 195.770000 81.800000 ;
      RECT 143.560000 80.720000 186.760000 81.800000 ;
      RECT 98.560000 80.720000 141.760000 81.800000 ;
      RECT 53.560000 80.720000 96.760000 81.800000 ;
      RECT 8.560000 80.720000 51.760000 81.800000 ;
      RECT 4.330000 80.720000 6.760000 81.800000 ;
      RECT 1.000000 80.720000 2.530000 81.400000 ;
      RECT 1.000000 80.420000 199.100000 80.720000 ;
      RECT 0.000000 80.180000 200.100000 80.420000 ;
      RECT 1.000000 79.200000 199.100000 80.180000 ;
      RECT 0.000000 79.080000 200.100000 79.200000 ;
      RECT 199.370000 78.350000 200.100000 79.080000 ;
      RECT 0.000000 78.350000 0.730000 79.080000 ;
      RECT 186.560000 78.000000 197.570000 79.080000 ;
      RECT 141.560000 78.000000 184.760000 79.080000 ;
      RECT 96.560000 78.000000 139.760000 79.080000 ;
      RECT 51.560000 78.000000 94.760000 79.080000 ;
      RECT 6.560000 78.000000 49.760000 79.080000 ;
      RECT 2.530000 78.000000 4.595000 79.080000 ;
      RECT 1.000000 77.370000 199.100000 78.000000 ;
      RECT 0.000000 77.130000 200.100000 77.370000 ;
      RECT 1.000000 76.360000 199.100000 77.130000 ;
      RECT 197.570000 76.150000 199.100000 76.360000 ;
      RECT 1.000000 76.150000 2.530000 76.360000 ;
      RECT 197.570000 75.300000 200.100000 76.150000 ;
      RECT 0.000000 75.300000 2.530000 76.150000 ;
      RECT 197.570000 75.280000 199.100000 75.300000 ;
      RECT 188.560000 75.280000 195.770000 76.360000 ;
      RECT 143.560000 75.280000 186.760000 76.360000 ;
      RECT 98.560000 75.280000 141.760000 76.360000 ;
      RECT 53.560000 75.280000 96.760000 76.360000 ;
      RECT 8.560000 75.280000 51.760000 76.360000 ;
      RECT 4.330000 75.280000 6.760000 76.360000 ;
      RECT 1.000000 75.280000 2.530000 75.300000 ;
      RECT 1.000000 74.320000 199.100000 75.280000 ;
      RECT 0.000000 74.080000 200.100000 74.320000 ;
      RECT 1.000000 73.640000 199.100000 74.080000 ;
      RECT 199.370000 72.560000 200.100000 73.100000 ;
      RECT 186.560000 72.560000 197.570000 73.640000 ;
      RECT 141.560000 72.560000 184.760000 73.640000 ;
      RECT 96.560000 72.560000 139.760000 73.640000 ;
      RECT 51.560000 72.560000 94.760000 73.640000 ;
      RECT 6.560000 72.560000 49.760000 73.640000 ;
      RECT 2.530000 72.560000 4.595000 73.640000 ;
      RECT 0.000000 72.560000 0.730000 73.100000 ;
      RECT 0.000000 72.250000 200.100000 72.560000 ;
      RECT 1.000000 71.270000 199.100000 72.250000 ;
      RECT 0.000000 71.030000 200.100000 71.270000 ;
      RECT 1.000000 70.920000 199.100000 71.030000 ;
      RECT 197.570000 70.050000 199.100000 70.920000 ;
      RECT 1.000000 70.050000 2.530000 70.920000 ;
      RECT 197.570000 69.840000 200.100000 70.050000 ;
      RECT 188.560000 69.840000 195.770000 70.920000 ;
      RECT 143.560000 69.840000 186.760000 70.920000 ;
      RECT 98.560000 69.840000 141.760000 70.920000 ;
      RECT 53.560000 69.840000 96.760000 70.920000 ;
      RECT 8.560000 69.840000 51.760000 70.920000 ;
      RECT 4.330000 69.840000 6.760000 70.920000 ;
      RECT 0.000000 69.840000 2.530000 70.050000 ;
      RECT 0.000000 69.200000 200.100000 69.840000 ;
      RECT 1.000000 68.220000 199.100000 69.200000 ;
      RECT 0.000000 68.200000 200.100000 68.220000 ;
      RECT 199.370000 67.980000 200.100000 68.200000 ;
      RECT 0.000000 67.980000 0.730000 68.200000 ;
      RECT 186.560000 67.120000 197.570000 68.200000 ;
      RECT 141.560000 67.120000 184.760000 68.200000 ;
      RECT 96.560000 67.120000 139.760000 68.200000 ;
      RECT 51.560000 67.120000 94.760000 68.200000 ;
      RECT 6.560000 67.120000 49.760000 68.200000 ;
      RECT 2.530000 67.120000 4.595000 68.200000 ;
      RECT 1.000000 67.000000 199.100000 67.120000 ;
      RECT 0.000000 66.760000 200.100000 67.000000 ;
      RECT 1.000000 65.780000 199.100000 66.760000 ;
      RECT 0.000000 65.480000 200.100000 65.780000 ;
      RECT 197.570000 64.930000 200.100000 65.480000 ;
      RECT 0.000000 64.930000 2.530000 65.480000 ;
      RECT 197.570000 64.400000 199.100000 64.930000 ;
      RECT 188.560000 64.400000 195.770000 65.480000 ;
      RECT 143.560000 64.400000 186.760000 65.480000 ;
      RECT 98.560000 64.400000 141.760000 65.480000 ;
      RECT 53.560000 64.400000 96.760000 65.480000 ;
      RECT 8.560000 64.400000 51.760000 65.480000 ;
      RECT 4.330000 64.400000 6.760000 65.480000 ;
      RECT 1.000000 64.400000 2.530000 64.930000 ;
      RECT 1.000000 63.950000 199.100000 64.400000 ;
      RECT 0.000000 63.710000 200.100000 63.950000 ;
      RECT 1.000000 62.760000 199.100000 63.710000 ;
      RECT 199.370000 61.880000 200.100000 62.730000 ;
      RECT 0.000000 61.880000 0.730000 62.730000 ;
      RECT 186.560000 61.680000 197.570000 62.760000 ;
      RECT 141.560000 61.680000 184.760000 62.760000 ;
      RECT 96.560000 61.680000 139.760000 62.760000 ;
      RECT 51.560000 61.680000 94.760000 62.760000 ;
      RECT 6.560000 61.680000 49.760000 62.760000 ;
      RECT 2.530000 61.680000 4.595000 62.760000 ;
      RECT 1.000000 60.900000 199.100000 61.680000 ;
      RECT 0.000000 60.660000 200.100000 60.900000 ;
      RECT 1.000000 60.040000 199.100000 60.660000 ;
      RECT 197.570000 59.680000 199.100000 60.040000 ;
      RECT 1.000000 59.680000 2.530000 60.040000 ;
      RECT 197.570000 58.960000 200.100000 59.680000 ;
      RECT 188.560000 58.960000 195.770000 60.040000 ;
      RECT 143.560000 58.960000 186.760000 60.040000 ;
      RECT 98.560000 58.960000 141.760000 60.040000 ;
      RECT 53.560000 58.960000 96.760000 60.040000 ;
      RECT 8.560000 58.960000 51.760000 60.040000 ;
      RECT 4.330000 58.960000 6.760000 60.040000 ;
      RECT 0.000000 58.960000 2.530000 59.680000 ;
      RECT 0.000000 58.830000 200.100000 58.960000 ;
      RECT 1.000000 57.850000 199.100000 58.830000 ;
      RECT 0.000000 57.610000 200.100000 57.850000 ;
      RECT 1.000000 57.320000 199.100000 57.610000 ;
      RECT 199.370000 56.240000 200.100000 56.630000 ;
      RECT 186.560000 56.240000 197.570000 57.320000 ;
      RECT 141.560000 56.240000 184.760000 57.320000 ;
      RECT 96.560000 56.240000 139.760000 57.320000 ;
      RECT 51.560000 56.240000 94.760000 57.320000 ;
      RECT 6.560000 56.240000 49.760000 57.320000 ;
      RECT 2.530000 56.240000 4.595000 57.320000 ;
      RECT 0.000000 56.240000 0.730000 56.630000 ;
      RECT 0.000000 55.780000 200.100000 56.240000 ;
      RECT 1.000000 54.800000 199.100000 55.780000 ;
      RECT 0.000000 54.600000 200.100000 54.800000 ;
      RECT 197.570000 54.560000 200.100000 54.600000 ;
      RECT 0.000000 54.560000 2.530000 54.600000 ;
      RECT 197.570000 53.580000 199.100000 54.560000 ;
      RECT 1.000000 53.580000 2.530000 54.560000 ;
      RECT 197.570000 53.520000 200.100000 53.580000 ;
      RECT 188.560000 53.520000 195.770000 54.600000 ;
      RECT 143.560000 53.520000 186.760000 54.600000 ;
      RECT 98.560000 53.520000 141.760000 54.600000 ;
      RECT 53.560000 53.520000 96.760000 54.600000 ;
      RECT 8.560000 53.520000 51.760000 54.600000 ;
      RECT 4.330000 53.520000 6.760000 54.600000 ;
      RECT 0.000000 53.520000 2.530000 53.580000 ;
      RECT 0.000000 53.340000 200.100000 53.520000 ;
      RECT 1.000000 52.360000 199.100000 53.340000 ;
      RECT 0.000000 51.880000 200.100000 52.360000 ;
      RECT 199.370000 51.510000 200.100000 51.880000 ;
      RECT 0.000000 51.510000 0.730000 51.880000 ;
      RECT 186.560000 50.800000 197.570000 51.880000 ;
      RECT 141.560000 50.800000 184.760000 51.880000 ;
      RECT 96.560000 50.800000 139.760000 51.880000 ;
      RECT 51.560000 50.800000 94.760000 51.880000 ;
      RECT 6.560000 50.800000 49.760000 51.880000 ;
      RECT 2.530000 50.800000 4.595000 51.880000 ;
      RECT 1.000000 50.530000 199.100000 50.800000 ;
      RECT 0.000000 50.290000 200.100000 50.530000 ;
      RECT 1.000000 49.310000 199.100000 50.290000 ;
      RECT 0.000000 49.160000 200.100000 49.310000 ;
      RECT 197.570000 48.460000 200.100000 49.160000 ;
      RECT 0.000000 48.460000 2.530000 49.160000 ;
      RECT 197.570000 48.080000 199.100000 48.460000 ;
      RECT 188.560000 48.080000 195.770000 49.160000 ;
      RECT 143.560000 48.080000 186.760000 49.160000 ;
      RECT 98.560000 48.080000 141.760000 49.160000 ;
      RECT 53.560000 48.080000 96.760000 49.160000 ;
      RECT 8.560000 48.080000 51.760000 49.160000 ;
      RECT 4.330000 48.080000 6.760000 49.160000 ;
      RECT 1.000000 48.080000 2.530000 48.460000 ;
      RECT 1.000000 47.480000 199.100000 48.080000 ;
      RECT 0.000000 47.240000 200.100000 47.480000 ;
      RECT 1.000000 46.440000 199.100000 47.240000 ;
      RECT 199.370000 45.410000 200.100000 46.260000 ;
      RECT 0.000000 45.410000 0.730000 46.260000 ;
      RECT 186.560000 45.360000 197.570000 46.440000 ;
      RECT 141.560000 45.360000 184.760000 46.440000 ;
      RECT 96.560000 45.360000 139.760000 46.440000 ;
      RECT 51.560000 45.360000 94.760000 46.440000 ;
      RECT 6.560000 45.360000 49.760000 46.440000 ;
      RECT 2.530000 45.360000 4.595000 46.440000 ;
      RECT 1.000000 44.430000 199.100000 45.360000 ;
      RECT 0.000000 44.190000 200.100000 44.430000 ;
      RECT 1.000000 43.720000 199.100000 44.190000 ;
      RECT 197.570000 43.210000 199.100000 43.720000 ;
      RECT 1.000000 43.210000 2.530000 43.720000 ;
      RECT 197.570000 42.970000 200.100000 43.210000 ;
      RECT 0.000000 42.970000 2.530000 43.210000 ;
      RECT 197.570000 42.640000 199.100000 42.970000 ;
      RECT 188.560000 42.640000 195.770000 43.720000 ;
      RECT 143.560000 42.640000 186.760000 43.720000 ;
      RECT 98.560000 42.640000 141.760000 43.720000 ;
      RECT 53.560000 42.640000 96.760000 43.720000 ;
      RECT 8.560000 42.640000 51.760000 43.720000 ;
      RECT 4.330000 42.640000 6.760000 43.720000 ;
      RECT 1.000000 42.640000 2.530000 42.970000 ;
      RECT 1.000000 41.990000 199.100000 42.640000 ;
      RECT 0.000000 41.140000 200.100000 41.990000 ;
      RECT 1.000000 41.000000 199.100000 41.140000 ;
      RECT 199.370000 39.920000 200.100000 40.160000 ;
      RECT 186.560000 39.920000 197.570000 41.000000 ;
      RECT 141.560000 39.920000 184.760000 41.000000 ;
      RECT 96.560000 39.920000 139.760000 41.000000 ;
      RECT 51.560000 39.920000 94.760000 41.000000 ;
      RECT 6.560000 39.920000 49.760000 41.000000 ;
      RECT 2.530000 39.920000 4.595000 41.000000 ;
      RECT 0.000000 39.920000 0.730000 40.160000 ;
      RECT 1.000000 38.940000 199.100000 39.920000 ;
      RECT 0.000000 38.280000 200.100000 38.940000 ;
      RECT 197.570000 38.090000 200.100000 38.280000 ;
      RECT 0.000000 38.090000 2.530000 38.280000 ;
      RECT 197.570000 37.200000 199.100000 38.090000 ;
      RECT 188.560000 37.200000 195.770000 38.280000 ;
      RECT 143.560000 37.200000 186.760000 38.280000 ;
      RECT 98.560000 37.200000 141.760000 38.280000 ;
      RECT 53.560000 37.200000 96.760000 38.280000 ;
      RECT 8.560000 37.200000 51.760000 38.280000 ;
      RECT 4.330000 37.200000 6.760000 38.280000 ;
      RECT 1.000000 37.200000 2.530000 38.090000 ;
      RECT 1.000000 37.110000 199.100000 37.200000 ;
      RECT 0.000000 36.870000 200.100000 37.110000 ;
      RECT 1.000000 35.890000 199.100000 36.870000 ;
      RECT 0.000000 35.560000 200.100000 35.890000 ;
      RECT 199.370000 35.040000 200.100000 35.560000 ;
      RECT 0.000000 35.040000 0.730000 35.560000 ;
      RECT 186.560000 34.480000 197.570000 35.560000 ;
      RECT 141.560000 34.480000 184.760000 35.560000 ;
      RECT 96.560000 34.480000 139.760000 35.560000 ;
      RECT 51.560000 34.480000 94.760000 35.560000 ;
      RECT 6.560000 34.480000 49.760000 35.560000 ;
      RECT 2.530000 34.480000 4.595000 35.560000 ;
      RECT 1.000000 34.060000 199.100000 34.480000 ;
      RECT 0.000000 33.820000 200.100000 34.060000 ;
      RECT 1.000000 32.840000 199.100000 33.820000 ;
      RECT 197.570000 31.990000 200.100000 32.840000 ;
      RECT 0.000000 31.990000 2.530000 32.840000 ;
      RECT 197.570000 31.760000 199.100000 31.990000 ;
      RECT 188.560000 31.760000 195.770000 32.840000 ;
      RECT 143.560000 31.760000 186.760000 32.840000 ;
      RECT 98.560000 31.760000 141.760000 32.840000 ;
      RECT 53.560000 31.760000 96.760000 32.840000 ;
      RECT 8.560000 31.760000 51.760000 32.840000 ;
      RECT 4.330000 31.760000 6.760000 32.840000 ;
      RECT 1.000000 31.760000 2.530000 31.990000 ;
      RECT 1.000000 31.010000 199.100000 31.760000 ;
      RECT 0.000000 30.770000 200.100000 31.010000 ;
      RECT 1.000000 30.120000 199.100000 30.770000 ;
      RECT 199.370000 29.550000 200.100000 29.790000 ;
      RECT 0.000000 29.550000 0.730000 29.790000 ;
      RECT 186.560000 29.040000 197.570000 30.120000 ;
      RECT 141.560000 29.040000 184.760000 30.120000 ;
      RECT 96.560000 29.040000 139.760000 30.120000 ;
      RECT 51.560000 29.040000 94.760000 30.120000 ;
      RECT 6.560000 29.040000 49.760000 30.120000 ;
      RECT 2.530000 29.040000 4.595000 30.120000 ;
      RECT 1.000000 28.570000 199.100000 29.040000 ;
      RECT 0.000000 27.720000 200.100000 28.570000 ;
      RECT 1.000000 27.400000 199.100000 27.720000 ;
      RECT 197.570000 26.740000 199.100000 27.400000 ;
      RECT 1.000000 26.740000 2.530000 27.400000 ;
      RECT 197.570000 26.500000 200.100000 26.740000 ;
      RECT 0.000000 26.500000 2.530000 26.740000 ;
      RECT 197.570000 26.320000 199.100000 26.500000 ;
      RECT 188.560000 26.320000 195.770000 27.400000 ;
      RECT 143.560000 26.320000 186.760000 27.400000 ;
      RECT 98.560000 26.320000 141.760000 27.400000 ;
      RECT 53.560000 26.320000 96.760000 27.400000 ;
      RECT 8.560000 26.320000 51.760000 27.400000 ;
      RECT 4.330000 26.320000 6.760000 27.400000 ;
      RECT 1.000000 26.320000 2.530000 26.500000 ;
      RECT 1.000000 25.520000 199.100000 26.320000 ;
      RECT 0.000000 24.680000 200.100000 25.520000 ;
      RECT 199.370000 24.670000 200.100000 24.680000 ;
      RECT 0.000000 24.670000 0.730000 24.680000 ;
      RECT 199.370000 23.600000 200.100000 23.690000 ;
      RECT 186.560000 23.600000 197.570000 24.680000 ;
      RECT 141.560000 23.600000 184.760000 24.680000 ;
      RECT 96.560000 23.600000 139.760000 24.680000 ;
      RECT 51.560000 23.600000 94.760000 24.680000 ;
      RECT 6.560000 23.600000 49.760000 24.680000 ;
      RECT 2.530000 23.600000 4.595000 24.680000 ;
      RECT 0.000000 23.600000 0.730000 23.690000 ;
      RECT 0.000000 23.450000 200.100000 23.600000 ;
      RECT 1.000000 22.470000 199.100000 23.450000 ;
      RECT 0.000000 21.960000 200.100000 22.470000 ;
      RECT 197.570000 21.620000 200.100000 21.960000 ;
      RECT 0.000000 21.620000 2.530000 21.960000 ;
      RECT 197.570000 20.880000 199.100000 21.620000 ;
      RECT 188.560000 20.880000 195.770000 21.960000 ;
      RECT 143.560000 20.880000 186.760000 21.960000 ;
      RECT 98.560000 20.880000 141.760000 21.960000 ;
      RECT 53.560000 20.880000 96.760000 21.960000 ;
      RECT 8.560000 20.880000 51.760000 21.960000 ;
      RECT 4.330000 20.880000 6.760000 21.960000 ;
      RECT 1.000000 20.880000 2.530000 21.620000 ;
      RECT 1.000000 20.640000 199.100000 20.880000 ;
      RECT 0.000000 20.400000 200.100000 20.640000 ;
      RECT 1.000000 19.420000 199.100000 20.400000 ;
      RECT 0.000000 19.240000 200.100000 19.420000 ;
      RECT 199.370000 18.570000 200.100000 19.240000 ;
      RECT 0.000000 18.570000 0.730000 19.240000 ;
      RECT 186.560000 18.160000 197.570000 19.240000 ;
      RECT 141.560000 18.160000 184.760000 19.240000 ;
      RECT 96.560000 18.160000 139.760000 19.240000 ;
      RECT 51.560000 18.160000 94.760000 19.240000 ;
      RECT 6.560000 18.160000 49.760000 19.240000 ;
      RECT 2.530000 18.160000 4.595000 19.240000 ;
      RECT 1.000000 17.590000 199.100000 18.160000 ;
      RECT 0.000000 17.350000 200.100000 17.590000 ;
      RECT 1.000000 16.520000 199.100000 17.350000 ;
      RECT 197.570000 16.370000 199.100000 16.520000 ;
      RECT 1.000000 16.370000 2.530000 16.520000 ;
      RECT 197.570000 16.130000 200.100000 16.370000 ;
      RECT 0.000000 16.130000 2.530000 16.370000 ;
      RECT 197.570000 15.440000 199.100000 16.130000 ;
      RECT 188.560000 15.440000 195.770000 16.520000 ;
      RECT 143.560000 15.440000 186.760000 16.520000 ;
      RECT 98.560000 15.440000 141.760000 16.520000 ;
      RECT 53.560000 15.440000 96.760000 16.520000 ;
      RECT 8.560000 15.440000 51.760000 16.520000 ;
      RECT 4.330000 15.440000 6.760000 16.520000 ;
      RECT 1.000000 15.440000 2.530000 16.130000 ;
      RECT 1.000000 15.150000 199.100000 15.440000 ;
      RECT 0.000000 14.300000 200.100000 15.150000 ;
      RECT 1.000000 13.800000 199.100000 14.300000 ;
      RECT 199.370000 13.080000 200.100000 13.320000 ;
      RECT 0.000000 13.080000 0.730000 13.320000 ;
      RECT 186.560000 12.720000 197.570000 13.800000 ;
      RECT 141.560000 12.720000 184.760000 13.800000 ;
      RECT 96.560000 12.720000 139.760000 13.800000 ;
      RECT 51.560000 12.720000 94.760000 13.800000 ;
      RECT 6.560000 12.720000 49.760000 13.800000 ;
      RECT 2.530000 12.720000 4.595000 13.800000 ;
      RECT 1.000000 12.100000 199.100000 12.720000 ;
      RECT 0.000000 11.250000 200.100000 12.100000 ;
      RECT 1.000000 11.080000 199.100000 11.250000 ;
      RECT 197.570000 10.270000 199.100000 11.080000 ;
      RECT 1.000000 10.270000 2.530000 11.080000 ;
      RECT 197.570000 10.030000 200.100000 10.270000 ;
      RECT 0.000000 10.030000 2.530000 10.270000 ;
      RECT 197.570000 10.000000 199.100000 10.030000 ;
      RECT 188.560000 10.000000 195.770000 11.080000 ;
      RECT 143.560000 10.000000 186.760000 11.080000 ;
      RECT 98.560000 10.000000 141.760000 11.080000 ;
      RECT 53.560000 10.000000 96.760000 11.080000 ;
      RECT 8.560000 10.000000 51.760000 11.080000 ;
      RECT 4.330000 10.000000 6.760000 11.080000 ;
      RECT 1.000000 10.000000 2.530000 10.030000 ;
      RECT 1.000000 9.050000 199.100000 10.000000 ;
      RECT 0.000000 8.360000 200.100000 9.050000 ;
      RECT 199.370000 8.200000 200.100000 8.360000 ;
      RECT 0.000000 8.200000 0.730000 8.360000 ;
      RECT 186.560000 7.280000 197.570000 8.360000 ;
      RECT 141.560000 7.280000 184.760000 8.360000 ;
      RECT 96.560000 7.280000 139.760000 8.360000 ;
      RECT 51.560000 7.280000 94.760000 8.360000 ;
      RECT 6.560000 7.280000 49.760000 8.360000 ;
      RECT 2.530000 7.280000 4.595000 8.360000 ;
      RECT 1.000000 7.220000 199.100000 7.280000 ;
      RECT 0.000000 6.980000 200.100000 7.220000 ;
      RECT 1.000000 6.000000 199.100000 6.980000 ;
      RECT 0.000000 5.760000 200.100000 6.000000 ;
      RECT 1.000000 5.640000 199.100000 5.760000 ;
      RECT 197.570000 4.780000 199.100000 5.640000 ;
      RECT 1.000000 4.780000 2.530000 5.640000 ;
      RECT 197.570000 4.560000 200.100000 4.780000 ;
      RECT 188.560000 4.560000 195.770000 5.640000 ;
      RECT 143.560000 4.560000 186.760000 5.640000 ;
      RECT 98.560000 4.560000 141.760000 5.640000 ;
      RECT 53.560000 4.560000 96.760000 5.640000 ;
      RECT 8.560000 4.560000 51.760000 5.640000 ;
      RECT 4.330000 4.560000 6.760000 5.640000 ;
      RECT 0.000000 4.560000 2.530000 4.780000 ;
      RECT 0.000000 4.350000 200.100000 4.560000 ;
      RECT 0.000000 0.000000 200.100000 0.750000 ;
    LAYER met4 ;
      RECT 4.330000 198.320000 195.770000 200.260000 ;
      RECT 186.560000 196.520000 195.770000 198.320000 ;
      RECT 141.560000 196.520000 184.760000 198.320000 ;
      RECT 96.560000 196.520000 139.760000 198.320000 ;
      RECT 51.560000 196.520000 94.760000 198.320000 ;
      RECT 6.560000 196.520000 49.760000 198.320000 ;
      RECT 4.330000 193.320000 4.760000 198.320000 ;
      RECT 4.330000 192.240000 4.595000 193.320000 ;
      RECT 4.330000 187.880000 4.760000 192.240000 ;
      RECT 4.330000 186.800000 4.595000 187.880000 ;
      RECT 4.330000 182.440000 4.760000 186.800000 ;
      RECT 4.330000 181.360000 4.595000 182.440000 ;
      RECT 4.330000 177.000000 4.760000 181.360000 ;
      RECT 4.330000 175.920000 4.595000 177.000000 ;
      RECT 4.330000 171.560000 4.760000 175.920000 ;
      RECT 4.330000 170.480000 4.595000 171.560000 ;
      RECT 4.330000 166.120000 4.760000 170.480000 ;
      RECT 4.330000 165.040000 4.595000 166.120000 ;
      RECT 4.330000 160.680000 4.760000 165.040000 ;
      RECT 4.330000 159.600000 4.595000 160.680000 ;
      RECT 4.330000 155.240000 4.760000 159.600000 ;
      RECT 4.330000 154.160000 4.595000 155.240000 ;
      RECT 4.330000 149.800000 4.760000 154.160000 ;
      RECT 4.330000 148.720000 4.595000 149.800000 ;
      RECT 4.330000 144.360000 4.760000 148.720000 ;
      RECT 4.330000 143.280000 4.595000 144.360000 ;
      RECT 4.330000 138.920000 4.760000 143.280000 ;
      RECT 4.330000 137.840000 4.595000 138.920000 ;
      RECT 4.330000 133.480000 4.760000 137.840000 ;
      RECT 4.330000 132.400000 4.595000 133.480000 ;
      RECT 4.330000 128.040000 4.760000 132.400000 ;
      RECT 4.330000 126.960000 4.595000 128.040000 ;
      RECT 4.330000 122.600000 4.760000 126.960000 ;
      RECT 4.330000 121.520000 4.595000 122.600000 ;
      RECT 4.330000 117.160000 4.760000 121.520000 ;
      RECT 4.330000 116.080000 4.595000 117.160000 ;
      RECT 4.330000 111.720000 4.760000 116.080000 ;
      RECT 4.330000 110.640000 4.595000 111.720000 ;
      RECT 4.330000 106.280000 4.760000 110.640000 ;
      RECT 4.330000 105.200000 4.595000 106.280000 ;
      RECT 4.330000 100.840000 4.760000 105.200000 ;
      RECT 4.330000 99.760000 4.595000 100.840000 ;
      RECT 4.330000 95.400000 4.760000 99.760000 ;
      RECT 4.330000 94.320000 4.595000 95.400000 ;
      RECT 4.330000 89.960000 4.760000 94.320000 ;
      RECT 4.330000 88.880000 4.595000 89.960000 ;
      RECT 4.330000 84.520000 4.760000 88.880000 ;
      RECT 4.330000 83.440000 4.595000 84.520000 ;
      RECT 4.330000 79.080000 4.760000 83.440000 ;
      RECT 4.330000 78.000000 4.595000 79.080000 ;
      RECT 4.330000 73.640000 4.760000 78.000000 ;
      RECT 4.330000 72.560000 4.595000 73.640000 ;
      RECT 4.330000 68.200000 4.760000 72.560000 ;
      RECT 4.330000 67.120000 4.595000 68.200000 ;
      RECT 4.330000 62.760000 4.760000 67.120000 ;
      RECT 4.330000 61.680000 4.595000 62.760000 ;
      RECT 4.330000 57.320000 4.760000 61.680000 ;
      RECT 4.330000 56.240000 4.595000 57.320000 ;
      RECT 4.330000 51.880000 4.760000 56.240000 ;
      RECT 4.330000 50.800000 4.595000 51.880000 ;
      RECT 4.330000 46.440000 4.760000 50.800000 ;
      RECT 4.330000 45.360000 4.595000 46.440000 ;
      RECT 4.330000 41.000000 4.760000 45.360000 ;
      RECT 4.330000 39.920000 4.595000 41.000000 ;
      RECT 4.330000 35.560000 4.760000 39.920000 ;
      RECT 4.330000 34.480000 4.595000 35.560000 ;
      RECT 4.330000 30.120000 4.760000 34.480000 ;
      RECT 4.330000 29.040000 4.595000 30.120000 ;
      RECT 4.330000 24.680000 4.760000 29.040000 ;
      RECT 4.330000 23.600000 4.595000 24.680000 ;
      RECT 4.330000 19.240000 4.760000 23.600000 ;
      RECT 4.330000 18.160000 4.595000 19.240000 ;
      RECT 4.330000 13.800000 4.760000 18.160000 ;
      RECT 4.330000 12.720000 4.595000 13.800000 ;
      RECT 4.330000 8.360000 4.760000 12.720000 ;
      RECT 4.330000 7.280000 4.595000 8.360000 ;
      RECT 188.560000 2.550000 195.770000 196.520000 ;
      RECT 186.560000 2.550000 186.760000 196.520000 ;
      RECT 143.560000 2.550000 184.760000 196.520000 ;
      RECT 141.560000 2.550000 141.760000 196.520000 ;
      RECT 98.560000 2.550000 139.760000 196.520000 ;
      RECT 96.560000 2.550000 96.760000 196.520000 ;
      RECT 53.560000 2.550000 94.760000 196.520000 ;
      RECT 51.560000 2.550000 51.760000 196.520000 ;
      RECT 8.560000 2.550000 49.760000 196.520000 ;
      RECT 6.560000 2.550000 6.760000 196.520000 ;
      RECT 186.560000 0.750000 195.770000 2.550000 ;
      RECT 141.560000 0.750000 184.760000 2.550000 ;
      RECT 96.560000 0.750000 139.760000 2.550000 ;
      RECT 51.560000 0.750000 94.760000 2.550000 ;
      RECT 6.560000 0.750000 49.760000 2.550000 ;
      RECT 4.330000 0.750000 4.760000 7.280000 ;
      RECT 199.370000 0.000000 200.100000 200.260000 ;
      RECT 4.330000 0.000000 195.770000 0.750000 ;
      RECT 0.000000 0.000000 0.730000 200.260000 ;
  END
END RegFile

END LIBRARY
