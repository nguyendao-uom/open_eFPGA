##
## LEF for PtnCells ;
## created by Innovus v19.11-s128_1 on Mon Dec  6 12:36:37 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO LUT4AB
  CLASS BLOCK ;
  SIZE 200.100000 BY 200.260000 ;
  FOREIGN LUT4AB 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.027 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 9.240000 199.560000 9.620000 200.260000 ;
    END
  END N1BEG[3]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.4842 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.313 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 7.860000 199.560000 8.240000 200.260000 ;
    END
  END N1BEG[2]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0814 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.299 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 6.480000 199.560000 6.860000 200.260000 ;
    END
  END N1BEG[1]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9428 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.606 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 199.560000 5.480000 200.260000 ;
    END
  END N1BEG[0]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.843 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.107 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 21.660000 199.560000 22.040000 200.260000 ;
    END
  END N2BEG[7]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6218 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.001 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 19.820000 199.560000 20.200000 200.260000 ;
    END
  END N2BEG[6]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.129 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.537 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 18.440000 199.560000 18.820000 200.260000 ;
    END
  END N2BEG[5]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.679 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.169 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 17.060000 199.560000 17.440000 200.260000 ;
    END
  END N2BEG[4]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1482 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.633 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 15.680000 199.560000 16.060000 200.260000 ;
    END
  END N2BEG[3]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4622 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.203 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 13.840000 199.560000 14.220000 200.260000 ;
    END
  END N2BEG[2]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.129 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.537 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 12.460000 199.560000 12.840000 200.260000 ;
    END
  END N2BEG[1]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.323 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 11.080000 199.560000 11.460000 200.260000 ;
    END
  END N2BEG[0]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 33.620000 199.560000 34.000000 200.260000 ;
    END
  END N2BEGb[7]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7434 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.491 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 32.240000 199.560000 32.620000 200.260000 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5766 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.775 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 30.860000 199.560000 31.240000 200.260000 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.427 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.909 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 29.020000 199.560000 29.400000 200.260000 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.49 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 27.640000 199.560000 28.020000 200.260000 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0194 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.989 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 26.260000 199.560000 26.640000 200.260000 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 24.420000 199.560000 24.800000 200.260000 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.441 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 23.040000 199.560000 23.420000 200.260000 ;
    END
  END N2BEGb[0]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3046 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.415 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 58.000000 199.560000 58.380000 200.260000 ;
    END
  END N4BEG[15]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.5388 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.468 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 56.620000 199.560000 57.000000 200.260000 ;
    END
  END N4BEG[14]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6597 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.16 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.6978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 84.192 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 54.780000 199.560000 55.160000 200.260000 ;
    END
  END N4BEG[13]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.825 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.899 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 53.400000 199.560000 53.780000 200.260000 ;
    END
  END N4BEG[12]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.4825 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.1865 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 52.020000 199.560000 52.400000 200.260000 ;
    END
  END N4BEG[11]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.0442 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.995 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 50.180000 199.560000 50.560000 200.260000 ;
    END
  END N4BEG[10]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.3234 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.509 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 48.800000 199.560000 49.180000 200.260000 ;
    END
  END N4BEG[9]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6046 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.915 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 47.420000 199.560000 47.800000 200.260000 ;
    END
  END N4BEG[8]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.4138 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.961 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 45.580000 199.560000 45.960000 200.260000 ;
    END
  END N4BEG[7]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.971 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.747 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 44.200000 199.560000 44.580000 200.260000 ;
    END
  END N4BEG[6]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.5593 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.6885 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 42.820000 199.560000 43.200000 200.260000 ;
    END
  END N4BEG[5]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6524 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.036 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 41.440000 199.560000 41.820000 200.260000 ;
    END
  END N4BEG[4]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7434 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.491 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 39.600000 199.560000 39.980000 200.260000 ;
    END
  END N4BEG[3]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6314 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.931 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 38.220000 199.560000 38.600000 200.260000 ;
    END
  END N4BEG[2]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9557 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6705 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 36.840000 199.560000 37.220000 200.260000 ;
    END
  END N4BEG[1]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.129 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.537 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 35.000000 199.560000 35.380000 200.260000 ;
    END
  END N4BEG[0]
  PIN NN4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.679 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.169 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 82.380000 199.560000 82.760000 200.260000 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.4893 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.2855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.9976 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.928 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 80.540000 199.560000 80.920000 200.260000 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.813 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 79.160000 199.560000 79.540000 200.260000 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.315 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.349 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 77.780000 199.560000 78.160000 200.260000 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1458 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.621 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 75.940000 199.560000 76.320000 200.260000 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.027 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 74.560000 199.560000 74.940000 200.260000 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.6378 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.081 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 73.180000 199.560000 73.560000 200.260000 ;
    END
  END NN4BEG[9]
  PIN NN4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.323 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 71.800000 199.560000 72.180000 200.260000 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3362 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 69.960000 199.560000 70.340000 200.260000 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.843 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.107 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 68.580000 199.560000 68.960000 200.260000 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0814 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.299 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 67.200000 199.560000 67.580000 200.260000 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2982 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.265 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 65.360000 199.560000 65.740000 200.260000 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5266 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.525 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 63.980000 199.560000 64.360000 200.260000 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.829 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.037 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 62.600000 199.560000 62.980000 200.260000 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2578 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.181 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 60.760000 199.560000 61.140000 200.260000 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.441 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 59.380000 199.560000 59.760000 200.260000 ;
    END
  END NN4BEG[0]
  PIN Co
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4622 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.203 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 164.260000 199.560000 164.640000 200.260000 ;
    END
  END Co
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6355 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7805 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 7.8553 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.6372 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 8.474 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 24.8516 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.0085 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 317.52 LAYER met4  ;
    ANTENNAGATEAREA 2.0247 LAYER met4  ;
    ANTENNAMAXAREACAR 90.06 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 472.289 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 9.240000 0.000000 9.620000 0.700000 ;
    END
  END N1END[3]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.2365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.5595 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 20.6045 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 83.9133 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.390645 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.3344 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.912 LAYER met3  ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 23.7058 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 101.068 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.627985 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 58.3527 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 314.032 LAYER met4  ;
    ANTENNAGATEAREA 2.0247 LAYER met4  ;
    ANTENNAMAXAREACAR 80.1695 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 408.921 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.09371 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 7.860000 0.000000 8.240000 0.700000 ;
    END
  END N1END[2]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.4731 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.9785 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 13.2344 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 47.4005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.926 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.072 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 19.9655 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 84.3731 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.5145 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 245.552 LAYER met4  ;
    ANTENNAGATEAREA 2.0247 LAYER met4  ;
    ANTENNAMAXAREACAR 95.0293 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 499.888 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 6.480000 0.000000 6.860000 0.700000 ;
    END
  END N1END[1]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1595 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6055 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 10.3241 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.9641 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.446 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.512 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 15.951 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 64.0476 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.6006 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 132.144 LAYER met4  ;
    ANTENNAGATEAREA 2.0247 LAYER met4  ;
    ANTENNAMAXAREACAR 43.8101 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 216.085 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.674423 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 0.000000 5.480000 0.700000 ;
    END
  END N1END[0]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1731 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.7045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 69.9765 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 376.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8132 LAYER met4  ;
    ANTENNAMAXAREACAR 89.5912 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 457.607 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 21.660000 0.000000 22.040000 0.700000 ;
    END
  END N2MID[7]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.8515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.6771 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 309.488 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6542 LAYER met4  ;
    ANTENNAMAXAREACAR 87.2564 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 447.944 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 19.820000 0.000000 20.200000 0.700000 ;
    END
  END N2MID[6]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3477 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.5775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.1733 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 215.664 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8132 LAYER met4  ;
    ANTENNAMAXAREACAR 84.7327 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 438.048 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.637736 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 18.440000 0.000000 18.820000 0.700000 ;
    END
  END N2MID[5]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9051 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.0105 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met2  ;
    ANTENNAMAXAREACAR 23.7589 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 108.463 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.659431 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 24.0923 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 110.865 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.712573 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.3956 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 184.384 LAYER met4  ;
    ANTENNAGATEAREA 1.6542 LAYER met4  ;
    ANTENNAMAXAREACAR 53.2199 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 276.879 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 17.060000 0.000000 17.440000 0.700000 ;
    END
  END N2MID[4]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.219 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.8358 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 74.1981 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.992 LAYER met3  ;
    ANTENNAGATEAREA 1.8132 LAYER met3  ;
    ANTENNAMAXAREACAR 17.5102 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 78.0543 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 15.680000 0.000000 16.060000 0.700000 ;
    END
  END N2MID[3]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.3295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 64.9263 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 347.68 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6542 LAYER met4  ;
    ANTENNAMAXAREACAR 76.2228 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 389.767 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.674423 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 13.840000 0.000000 14.220000 0.700000 ;
    END
  END N2MID[2]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.6407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.1285 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0707 LAYER met2  ;
    ANTENNAMAXAREACAR 12.0276 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 50.1831 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.360629 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAGATEAREA 1.0707 LAYER met3  ;
    ANTENNAMAXAREACAR 12.4012 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 52.6114 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.397988 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.0246 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 273.072 LAYER met4  ;
    ANTENNAGATEAREA 1.8132 LAYER met4  ;
    ANTENNAMAXAREACAR 40.5418 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 203.214 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.397988 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 12.460000 0.000000 12.840000 0.700000 ;
    END
  END N2MID[1]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.9362 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.229 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6542 LAYER met2  ;
    ANTENNAMAXAREACAR 12.6896 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 54.9168 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 11.080000 0.000000 11.460000 0.700000 ;
    END
  END N2MID[0]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1327 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.1585 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 11.2995 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.6098 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 11.9182 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 41.8242 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 58.3308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 313.44 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 79.9555 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 421.707 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 33.620000 0.000000 34.000000 0.700000 ;
    END
  END N2END[7]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5203 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3325 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 8.29768 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.9883 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.263 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.536 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 13.5036 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 51.8265 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.9064 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 192.912 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 87.326 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 440.777 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.857862 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 32.240000 0.000000 32.620000 0.700000 ;
    END
  END N2END[6]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2947 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.1945 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 13.9827 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 51.2974 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.492 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.424 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 31.2176 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 144.29 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.5717 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 232.848 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 66.6504 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 333.644 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 30.860000 0.000000 31.240000 0.700000 ;
    END
  END N2END[5]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.6615 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.3505 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met2  ;
    ANTENNAMAXAREACAR 22.1197 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 101.276 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.497308 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAGATEAREA 1.3887 LAYER met3  ;
    ANTENNAMAXAREACAR 22.6027 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 104.191 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 29.020000 0.000000 29.400000 0.700000 ;
    END
  END N2END[4]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 8.14125 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.1831 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2415 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.576 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 8.6968 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 25.8086 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.5448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 195.376 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 50.6434 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 252.727 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.548637 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 27.640000 0.000000 28.020000 0.700000 ;
    END
  END N2END[3]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.0383 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 79.0965 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0707 LAYER met2  ;
    ANTENNAMAXAREACAR 25.261 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 117.525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.502139 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.0508 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.408 LAYER met3  ;
    ANTENNAGATEAREA 1.2297 LAYER met3  ;
    ANTENNAMAXAREACAR 26.9288 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 126.802 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 26.260000 0.000000 26.640000 0.700000 ;
    END
  END N2END[2]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7807 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.1725 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met2  ;
    ANTENNAMAXAREACAR 37.2475 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 176.86 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.449057 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.87892 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.48 LAYER met3  ;
    ANTENNAGATEAREA 0.318 LAYER met3  ;
    ANTENNAMAXAREACAR 43.1561 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 209.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 43.6991 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 213.095 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 24.420000 0.000000 24.800000 0.700000 ;
    END
  END N2END[1]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 17.1797 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 85.0395 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met2  ;
    ANTENNAMAXAREACAR 43.3014 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 207.807 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.508654 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.5609 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.12 LAYER met3  ;
    ANTENNAGATEAREA 1.0707 LAYER met3  ;
    ANTENNAMAXAREACAR 48.4952 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 235.938 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.612202 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 71.4118 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 361.124 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 23.040000 0.000000 23.420000 0.700000 ;
    END
  END N2END[0]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6057 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7595 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 8.19784 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.4891 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.472 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 17.6894 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 74.1845 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.3176 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 103.968 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 36.5433 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 188.389 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 58.000000 0.000000 58.380000 0.700000 ;
    END
  END N4END[15]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9593 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4905 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 6.71083 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.9689 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 7.47228 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 20.1035 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.1478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 246.592 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 46.6736 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 233.298 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 56.620000 0.000000 57.000000 0.700000 ;
    END
  END N4END[14]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5031 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.2465 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 11.5956 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.4778 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 12.357 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 44.6124 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.9278 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 234.752 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 49.6725 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 244.028 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 54.780000 0.000000 55.160000 0.700000 ;
    END
  END N4END[13]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3743 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.6025 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 11.2993 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.9963 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.335725 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.256 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 12.0716 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 43.1861 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.9266 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 267.216 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 54.4829 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 270.179 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 53.400000 0.000000 53.780000 0.700000 ;
    END
  END N4END[12]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.5227 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.2165 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 12.6961 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.4375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 13.9337 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 52.1118 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.0608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 214.128 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 47.9643 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 234.008 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 52.020000 0.000000 52.400000 0.700000 ;
    END
  END N4END[11]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4222 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.767 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 14.2865 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 53.0806 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.236485 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 50.180000 0.000000 50.560000 0.700000 ;
    END
  END N4END[10]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.5441 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 117.387 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 25.6893 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 110.281 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.118242 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 48.800000 0.000000 49.180000 0.700000 ;
    END
  END N4END[9]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8275 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.8685 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 14.0497 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 51.7483 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 15.9222 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 62.8088 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.8046 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 261.232 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 57.3805 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 284.718 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 47.420000 0.000000 47.800000 0.700000 ;
    END
  END N4END[8]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6079 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6525 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 11.2441 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.4488 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 11.8307 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 41.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.5126 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 265.008 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 53.8903 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 266.725 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 45.580000 0.000000 45.960000 0.700000 ;
    END
  END N4END[7]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9135 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 9.00943 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.547 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 10.2471 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 34.2213 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.2848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 284.656 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 55.5111 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 276.029 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 44.200000 0.000000 44.580000 0.700000 ;
    END
  END N4END[6]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4165 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 8.98321 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.1445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 9.90338 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 32.1256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 55.7598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 297.856 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 57.2698 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 285.146 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 42.820000 0.000000 43.200000 0.700000 ;
    END
  END N4END[5]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2931 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.1965 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 10.668 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.8401 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.056 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.432 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 15.3977 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 61.1387 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.6618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 276 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 59.2831 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 295.593 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 41.440000 0.000000 41.820000 0.700000 ;
    END
  END N4END[4]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.9063 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.1345 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 13.0791 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.7564 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 13.6657 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 50.9156 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.7604 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 186.8 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 49.0337 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 249.539 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 39.600000 0.000000 39.980000 0.700000 ;
    END
  END N4END[3]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.6175 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.8185 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 17.6375 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 69.6871 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 19.3513 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 79.9011 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.679 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 192.16 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 116.24 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 611.731 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 38.220000 0.000000 38.600000 0.700000 ;
    END
  END N4END[2]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.505 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 81.011 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met2  ;
    ANTENNAMAXAREACAR 27.6688 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 129.998 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.606289 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 36.840000 0.000000 37.220000 0.700000 ;
    END
  END N4END[1]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.5477 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.8895 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met2  ;
    ANTENNAMAXAREACAR 15.5642 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 70.4025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.508654 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 27.4239 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 146.704 LAYER met3  ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 45.6442 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 231.315 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.552528 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 46.0385 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 233.8 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 35.000000 0.000000 35.380000 0.700000 ;
    END
  END N4END[0]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.2629 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.9275 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 20.8008 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 85.3876 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 23.6257 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 101.527 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.6078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 195.712 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 54.7231 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 267.78 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 82.380000 0.000000 82.760000 0.700000 ;
    END
  END NN4END[15]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.4939 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.2005 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 14.4309 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 53.8095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 17.5733 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 71.6425 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.0758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 262.208 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 59.2619 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 294.381 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 80.540000 0.000000 80.920000 0.700000 ;
    END
  END NN4END[14]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.3195 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.3185 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 14.7702 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 55.2346 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 15.3474 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 59.3938 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.2898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 194.016 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 46.1746 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 224.205 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 79.160000 0.000000 79.540000 0.700000 ;
    END
  END NN4END[13]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.3845 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 76.6535 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 39.484 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 179.075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 40.8804 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 187.596 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.2748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 129.936 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 61.5012 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 297.973 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 77.780000 0.000000 78.160000 0.700000 ;
    END
  END NN4END[12]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5245 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3535 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 8.30734 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.0366 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.24 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 17.2675 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 71.8979 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.1978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 300.192 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 65.0061 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 326.903 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 75.940000 0.000000 76.320000 0.700000 ;
    END
  END NN4END[11]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5245 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3535 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 9.64067 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.7032 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 10.7196 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 36.5309 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.2848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 284.656 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 55.9836 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 278.339 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 74.560000 0.000000 74.940000 0.700000 ;
    END
  END NN4END[10]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9493 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4675 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 9.52588 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 28.8578 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 10.1125 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 33.017 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 54.2238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 289.664 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 56.1742 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 279.079 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 73.180000 0.000000 73.560000 0.700000 ;
    END
  END NN4END[9]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2759 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.1105 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 11.8919 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.9593 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 14.8755 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 57.9457 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.0518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 278.08 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 59.0922 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 294.167 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 71.800000 0.000000 72.180000 0.700000 ;
    END
  END NN4END[8]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5675 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.5685 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 11.1511 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.2556 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.963 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.936 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 15.6669 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 62.4132 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.3536 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 264.16 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 57.5915 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 286.81 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 69.960000 0.000000 70.340000 0.700000 ;
    END
  END NN4END[7]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.395 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.706 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 8.30573 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.0285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.056 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 15.8926 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 64.5652 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.8688 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 261.104 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 57.4053 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 286.366 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 68.580000 0.000000 68.960000 0.700000 ;
    END
  END NN4END[6]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4866 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.207 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 28.7752 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 125.709 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.170002 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 67.200000 0.000000 67.580000 0.700000 ;
    END
  END NN4END[5]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.4691 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.0765 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 14.4104 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 53.5519 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 14.997 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 57.7111 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.0148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 267.216 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 57.4832 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 284.704 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 65.360000 0.000000 65.740000 0.700000 ;
    END
  END NN4END[4]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 18.1489 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 89.7575 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met2  ;
    ANTENNAMAXAREACAR 30.9803 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 144.622 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.517922 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.7038 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.224 LAYER met3  ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 35.0428 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 166.804 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 63.980000 0.000000 64.360000 0.700000 ;
    END
  END NN4END[3]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.8118 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 78.253 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met2  ;
    ANTENNAMAXAREACAR 26.2501 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 121.398 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.46478 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 62.600000 0.000000 62.980000 0.700000 ;
    END
  END NN4END[2]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.9069 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.1475 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 18.8326 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 75.5368 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.390645 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.067 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.824 LAYER met3  ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 23.9985 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 103.874 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.458019 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.7955 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 154.512 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 97.9769 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 507.999 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 60.760000 0.000000 61.140000 0.700000 ;
    END
  END NN4END[1]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.3754 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 81.179 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met2  ;
    ANTENNAMAXAREACAR 59.001 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 285.695 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.46478 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 59.380000 0.000000 59.760000 0.700000 ;
    END
  END NN4END[0]
  PIN Ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.7026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.179 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8082 LAYER met2  ;
    ANTENNAMAXAREACAR 11.4583 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.1003 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 164.260000 0.000000 164.640000 0.700000 ;
    END
  END Ci
  PIN E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 80.720000 200.100000 81.100000 ;
    END
  END E1BEG[3]
  PIN E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 79.500000 200.100000 79.880000 ;
    END
  END E1BEG[2]
  PIN E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 77.670000 200.100000 78.050000 ;
    END
  END E1BEG[1]
  PIN E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.3374 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 76.450000 200.100000 76.830000 ;
    END
  END E1BEG[0]
  PIN E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 92.920000 200.100000 93.300000 ;
    END
  END E2BEG[7]
  PIN E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.7914 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.216 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 91.090000 200.100000 91.470000 ;
    END
  END E2BEG[6]
  PIN E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 89.870000 200.100000 90.250000 ;
    END
  END E2BEG[5]
  PIN E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 88.040000 200.100000 88.420000 ;
    END
  END E2BEG[4]
  PIN E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 86.820000 200.100000 87.200000 ;
    END
  END E2BEG[3]
  PIN E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.8164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.016 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 84.990000 200.100000 85.370000 ;
    END
  END E2BEG[2]
  PIN E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 83.770000 200.100000 84.150000 ;
    END
  END E2BEG[1]
  PIN E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 81.940000 200.100000 82.320000 ;
    END
  END E2BEG[0]
  PIN E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 104.510000 200.100000 104.890000 ;
    END
  END E2BEGb[7]
  PIN E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 103.290000 200.100000 103.670000 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.656 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 101.460000 200.100000 101.840000 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 100.240000 200.100000 100.620000 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.2304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.224 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 98.410000 200.100000 98.790000 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 97.190000 200.100000 97.570000 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 95.360000 200.100000 95.740000 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.808 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 94.140000 200.100000 94.520000 ;
    END
  END E2BEGb[0]
  PIN EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.9064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.496 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 128.300000 200.100000 128.680000 ;
    END
  END EE4BEG[15]
  PIN EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.4138 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 127.080000 200.100000 127.460000 ;
    END
  END EE4BEG[14]
  PIN EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.4354 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.984 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 125.250000 200.100000 125.630000 ;
    END
  END EE4BEG[13]
  PIN EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5906 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 124.030000 200.100000 124.410000 ;
    END
  END EE4BEG[12]
  PIN EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 122.200000 200.100000 122.580000 ;
    END
  END EE4BEG[11]
  PIN EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.3314 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.096 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 120.980000 200.100000 121.360000 ;
    END
  END EE4BEG[10]
  PIN EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 119.150000 200.100000 119.530000 ;
    END
  END EE4BEG[9]
  PIN EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.656 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 117.930000 200.100000 118.310000 ;
    END
  END EE4BEG[8]
  PIN EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 116.710000 200.100000 117.090000 ;
    END
  END EE4BEG[7]
  PIN EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 114.880000 200.100000 115.260000 ;
    END
  END EE4BEG[6]
  PIN EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 113.660000 200.100000 114.040000 ;
    END
  END EE4BEG[5]
  PIN EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 111.830000 200.100000 112.210000 ;
    END
  END EE4BEG[4]
  PIN EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 110.610000 200.100000 110.990000 ;
    END
  END EE4BEG[3]
  PIN EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 108.780000 200.100000 109.160000 ;
    END
  END EE4BEG[2]
  PIN EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 107.560000 200.100000 107.940000 ;
    END
  END EE4BEG[1]
  PIN EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.1264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.336 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 105.730000 200.100000 106.110000 ;
    END
  END EE4BEG[0]
  PIN E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 145.990000 200.100000 146.370000 ;
    END
  END E6BEG[11]
  PIN E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 144.770000 200.100000 145.150000 ;
    END
  END E6BEG[10]
  PIN E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 143.550000 200.100000 143.930000 ;
    END
  END E6BEG[9]
  PIN E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.656 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 141.720000 200.100000 142.100000 ;
    END
  END E6BEG[8]
  PIN E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.0554 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.624 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 140.500000 200.100000 140.880000 ;
    END
  END E6BEG[7]
  PIN E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 138.670000 200.100000 139.050000 ;
    END
  END E6BEG[6]
  PIN E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.656 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 137.450000 200.100000 137.830000 ;
    END
  END E6BEG[5]
  PIN E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 135.620000 200.100000 136.000000 ;
    END
  END E6BEG[4]
  PIN E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.8384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.8 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 134.400000 200.100000 134.780000 ;
    END
  END E6BEG[3]
  PIN E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.1264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.336 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 132.570000 200.100000 132.950000 ;
    END
  END E6BEG[2]
  PIN E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 131.350000 200.100000 131.730000 ;
    END
  END E6BEG[1]
  PIN E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 130.130000 200.100000 130.510000 ;
    END
  END E6BEG[0]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4234 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.7399 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 192.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1837 LAYER met4  ;
    ANTENNAMAXAREACAR 81.6455 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 419.993 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 80.720000 0.700000 81.100000 ;
    END
  END E1END[3]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6816 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.2123 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 247.872 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1837 LAYER met4  ;
    ANTENNAMAXAREACAR 73.9504 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 379.906 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 79.500000 0.700000 79.880000 ;
    END
  END E1END[2]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 65.7117 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 353.28 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8657 LAYER met4  ;
    ANTENNAMAXAREACAR 114.993 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 607.909 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 77.670000 0.700000 78.050000 ;
    END
  END E1END[1]
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.2726 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.9106 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.464 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8657 LAYER met4  ;
    ANTENNAMAXAREACAR 36.153 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 179.265 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.744391 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 76.450000 0.700000 76.830000 ;
    END
  END E1END[0]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 33.5973 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 179.176 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8132 LAYER met3  ;
    ANTENNAMAXAREACAR 34.8168 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 171.874 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.493797 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 92.920000 0.700000 93.300000 ;
    END
  END E2MID[7]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.7884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 35.1702 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 163.954 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.512537 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.9356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 93.616 LAYER met4  ;
    ANTENNAGATEAREA 1.6542 LAYER met4  ;
    ANTENNAMAXAREACAR 60.9348 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 319.851 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 91.090000 0.700000 91.470000 ;
    END
  END E2MID[6]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 33.5838 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 180.032 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 64.397 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 328.905 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.769494 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.5415 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.824 LAYER met4  ;
    ANTENNAGATEAREA 1.8132 LAYER met4  ;
    ANTENNAMAXAREACAR 66.3502 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 339.838 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.769494 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 89.870000 0.700000 90.250000 ;
    END
  END E2MID[5]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.3825 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.36 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 24.8459 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 111.585 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 58.1382 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 313.824 LAYER met4  ;
    ANTENNAGATEAREA 1.6542 LAYER met4  ;
    ANTENNAMAXAREACAR 74.0326 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 392.658 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 88.040000 0.700000 88.420000 ;
    END
  END E2MID[4]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 55.162 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 294.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 75.248 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 398.723 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.1638 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 113.344 LAYER met4  ;
    ANTENNAGATEAREA 1.8132 LAYER met4  ;
    ANTENNAMAXAREACAR 86.9201 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 461.234 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.539497 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 86.820000 0.700000 87.200000 ;
    END
  END E2MID[3]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.8764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.136 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 57.2866 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 282.57 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    ANTENNAGATEAREA 1.6542 LAYER met4  ;
    ANTENNAMAXAREACAR 58.0222 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 286.777 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.481857 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 84.990000 0.700000 85.370000 ;
    END
  END E2MID[2]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.86 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.7246 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 159.472 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8132 LAYER met4  ;
    ANTENNAMAXAREACAR 50.4814 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 254.093 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.806793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 83.770000 0.700000 84.150000 ;
    END
  END E2MID[1]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0196 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.2621 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 152.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6542 LAYER met4  ;
    ANTENNAMAXAREACAR 52.6766 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 263.425 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.80021 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 81.940000 0.700000 82.320000 ;
    END
  END E2MID[0]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.5062 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.832 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met3  ;
    ANTENNAMAXAREACAR 39.1959 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 193.214 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.571064 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 104.510000 0.700000 104.890000 ;
    END
  END E2END[7]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.5568 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.44 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met3  ;
    ANTENNAMAXAREACAR 34.959 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 168.041 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 103.290000 0.700000 103.670000 ;
    END
  END E2END[6]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.503 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.952 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met3  ;
    ANTENNAMAXAREACAR 37.7341 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 185.53 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 101.460000 0.700000 101.840000 ;
    END
  END E2END[5]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.5338 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.984 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met3  ;
    ANTENNAMAXAREACAR 22.6421 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 109.496 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.515094 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 100.240000 0.700000 100.620000 ;
    END
  END E2END[4]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.2052 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 135.36 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 75.164 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 385.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.893789 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.4695 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.44 LAYER met4  ;
    ANTENNAGATEAREA 1.5477 LAYER met4  ;
    ANTENNAMAXAREACAR 79.3441 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 408.018 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.893789 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 98.410000 0.700000 98.790000 ;
    END
  END E2END[3]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8014 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.736 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 11.8799 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 42.0152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.5894 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.888 LAYER met4  ;
    ANTENNAGATEAREA 1.5477 LAYER met4  ;
    ANTENNAMAXAREACAR 38.2065 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 193.65 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 97.190000 0.700000 97.570000 ;
    END
  END E2END[2]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8906 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.3275 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 104.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0707 LAYER met4  ;
    ANTENNAMAXAREACAR 46.6255 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 233.548 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 95.360000 0.700000 95.740000 ;
    END
  END E2END[1]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0707 LAYER met3  ;
    ANTENNAMAXAREACAR 36.9092 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 178.984 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.527673 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 94.140000 0.700000 94.520000 ;
    END
  END E2END[0]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 40.4305 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 215.616 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 98.012 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 502.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.5958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.648 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 101.066 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 519.603 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 128.300000 0.700000 128.680000 ;
    END
  END EE4END[15]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 24.34 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 130.28 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 67.9324 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 340.483 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.6218 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 41.12 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 74.4069 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 375.413 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 127.080000 0.700000 127.460000 ;
    END
  END EE4END[14]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.8374 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.928 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 17.6273 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 73.2252 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.1646 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 183.152 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 46.6492 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 228.808 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 125.250000 0.700000 125.630000 ;
    END
  END EE4END[13]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 53.1192 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 283.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 52.7484 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 260.145 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 124.030000 0.700000 124.410000 ;
    END
  END EE4END[12]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 55.4538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 296.224 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 55.568 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 275.025 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 122.200000 0.700000 122.580000 ;
    END
  END EE4END[11]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 56.7972 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 303.384 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 54.8964 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 271.913 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 120.980000 0.700000 121.360000 ;
    END
  END EE4END[10]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 55.3692 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 295.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 57.6592 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 285.524 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.42052 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 119.150000 0.700000 119.530000 ;
    END
  END EE4END[9]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.9394 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.472 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 65.8208 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 311.655 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.5038 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 93.824 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 80.6898 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 391.356 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 117.930000 0.700000 118.310000 ;
    END
  END EE4END[8]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 54.2088 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 289.584 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 54.5576 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 269.691 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.42052 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 116.710000 0.700000 117.090000 ;
    END
  END EE4END[7]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 55.0932 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 294.296 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 60.4683 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 299.491 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.42052 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 114.880000 0.700000 115.260000 ;
    END
  END EE4END[6]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 32.9044 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 175.952 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 84.0147 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 427.723 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.1318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 85.8256 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 437.78 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 113.660000 0.700000 114.040000 ;
    END
  END EE4END[5]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 52.9188 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 282.704 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 58.4505 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 288.79 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.42052 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 111.830000 0.700000 112.210000 ;
    END
  END EE4END[4]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 95.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 67.2917 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 334.35 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 110.610000 0.700000 110.990000 ;
    END
  END EE4END[3]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.8722 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 111.784 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 65.9613 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 330.186 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.548637 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 108.780000 0.700000 109.160000 ;
    END
  END EE4END[2]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 55.4531 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 271.164 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.508654 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 107.560000 0.700000 107.940000 ;
    END
  END EE4END[1]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.3362 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 92.912 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 44.166 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 220.954 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.627985 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.0988 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 59.664 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 83.658 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 434.175 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 105.730000 0.700000 106.110000 ;
    END
  END EE4END[0]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 32.3554 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 173.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 83.3665 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 423.789 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.016 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 84.8119 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 432.297 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 145.990000 0.700000 146.370000 ;
    END
  END E6END[11]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 24.4672 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.424 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 64.4 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 324.274 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.512537 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.4978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.792 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 66.5219 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 335.99 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.512537 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 144.770000 0.700000 145.150000 ;
    END
  END E6END[10]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 44.2572 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 236.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 46.1078 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 231.404 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 143.550000 0.700000 143.930000 ;
    END
  END E6END[9]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.2135 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.792 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 37.193 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 178.583 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 55.6242 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 295.366 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 141.720000 0.700000 142.100000 ;
    END
  END E6END[8]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 57.2853 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 305.512 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 54.6412 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 271.144 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 140.500000 0.700000 140.880000 ;
    END
  END E6END[7]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 42.9899 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 213.377 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.152221 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 138.670000 0.700000 139.050000 ;
    END
  END E6END[6]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 53.6262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 286.472 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 53.3203 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 263.537 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 137.450000 0.700000 137.830000 ;
    END
  END E6END[5]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.877 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.144 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 48.5958 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 237.311 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.2506 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.944 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 50.5076 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 248.306 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 135.620000 0.700000 136.000000 ;
    END
  END E6END[4]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2514 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.136 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 16.4707 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 68.0308 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.5714 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 137.792 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 38.1929 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 185.081 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 134.400000 0.700000 134.780000 ;
    END
  END E6END[3]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 50.9928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 272.432 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 52.2639 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 257.069 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 132.570000 0.700000 132.950000 ;
    END
  END E6END[2]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 18.6743 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 76.5332 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.6611 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.736 LAYER met4  ;
    ANTENNAGATEAREA 2.3427 LAYER met4  ;
    ANTENNAMAXAREACAR 58.6842 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 304.987 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 131.350000 0.700000 131.730000 ;
    END
  END E6END[1]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.7254 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 15.0288 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 62.7306 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.666902 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.8927 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 106.56 LAYER met4  ;
    ANTENNAGATEAREA 2.3427 LAYER met4  ;
    ANTENNAMAXAREACAR 49.6179 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 244.73 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.666902 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 130.130000 0.700000 130.510000 ;
    END
  END E6END[0]
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.907 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 88.360000 0.000000 88.740000 0.700000 ;
    END
  END S1BEG[3]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1157 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4705 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 86.520000 0.000000 86.900000 0.700000 ;
    END
  END S1BEG[2]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.7506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.645 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 85.140000 0.000000 85.520000 0.700000 ;
    END
  END S1BEG[1]
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0602 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.075 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 83.760000 0.000000 84.140000 0.700000 ;
    END
  END S1BEG[0]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.344 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 112.740000 0.000000 113.120000 0.700000 ;
    END
  END S2BEG[7]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9174 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.361 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 110.900000 0.000000 111.280000 0.700000 ;
    END
  END S2BEG[6]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.599 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 109.520000 0.000000 109.900000 0.700000 ;
    END
  END S2BEG[5]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0674 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.229 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 108.140000 0.000000 108.520000 0.700000 ;
    END
  END S2BEG[4]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3794 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 106.300000 0.000000 106.680000 0.700000 ;
    END
  END S2BEG[3]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.621 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.997 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 104.920000 0.000000 105.300000 0.700000 ;
    END
  END S2BEG[2]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4102 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 103.540000 0.000000 103.920000 0.700000 ;
    END
  END S2BEG[1]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.871 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 101.700000 0.000000 102.080000 0.700000 ;
    END
  END S2BEG[0]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.189 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.719 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 100.320000 0.000000 100.700000 0.700000 ;
    END
  END S2BEGb[7]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8626 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.205 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 98.940000 0.000000 99.320000 0.700000 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7338 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.561 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 97.560000 0.000000 97.940000 0.700000 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4954 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.369 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 95.720000 0.000000 96.100000 0.700000 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3458 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.503 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 94.340000 0.000000 94.720000 0.700000 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.907 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 92.960000 0.000000 93.340000 0.700000 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.441 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 91.120000 0.000000 91.500000 0.700000 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3054 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.419 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 89.740000 0.000000 90.120000 0.700000 ;
    END
  END S2BEGb[0]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.8123 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.9535 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 136.660000 0.000000 137.040000 0.700000 ;
    END
  END S4BEG[15]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.6738 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.261 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 135.280000 0.000000 135.660000 0.700000 ;
    END
  END S4BEG[14]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.919 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.369 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 133.900000 0.000000 134.280000 0.700000 ;
    END
  END S4BEG[13]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.315 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.349 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 132.060000 0.000000 132.440000 0.700000 ;
    END
  END S4BEG[12]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.907 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 130.680000 0.000000 131.060000 0.700000 ;
    END
  END S4BEG[11]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.085 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 129.300000 0.000000 129.680000 0.700000 ;
    END
  END S4BEG[10]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 127.460000 0.000000 127.840000 0.700000 ;
    END
  END S4BEG[9]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3362 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 126.080000 0.000000 126.460000 0.700000 ;
    END
  END S4BEG[8]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.943 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.607 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 124.700000 0.000000 125.080000 0.700000 ;
    END
  END S4BEG[7]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.286 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 123.320000 0.000000 123.700000 0.700000 ;
    END
  END S4BEG[6]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0602 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.075 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 121.480000 0.000000 121.860000 0.700000 ;
    END
  END S4BEG[5]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6694 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.239 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 120.100000 0.000000 120.480000 0.700000 ;
    END
  END S4BEG[4]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.5139 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.4615 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 118.720000 0.000000 119.100000 0.700000 ;
    END
  END S4BEG[3]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1318 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.551 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 116.880000 0.000000 117.260000 0.700000 ;
    END
  END S4BEG[2]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.298 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 115.500000 0.000000 115.880000 0.700000 ;
    END
  END S4BEG[1]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.585 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 114.120000 0.000000 114.500000 0.700000 ;
    END
  END S4BEG[0]
  PIN SS4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.467 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 161.040000 0.000000 161.420000 0.700000 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.585 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 159.660000 0.000000 160.040000 0.700000 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1102 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.325 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.820000 0.000000 158.200000 0.700000 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.145 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 156.440000 0.000000 156.820000 0.700000 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.251 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 155.060000 0.000000 155.440000 0.700000 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.1474 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.629 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 153.680000 0.000000 154.060000 0.700000 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1766 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.775 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 151.840000 0.000000 152.220000 0.700000 ;
    END
  END SS4BEG[9]
  PIN SS4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6382 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.083 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.460000 0.000000 150.840000 0.700000 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.837 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 149.080000 0.000000 149.460000 0.700000 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2262 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.023 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 147.240000 0.000000 147.620000 0.700000 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.837 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 145.860000 0.000000 146.240000 0.700000 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.774 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 144.480000 0.000000 144.860000 0.700000 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4102 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 142.640000 0.000000 143.020000 0.700000 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7305 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.332 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.3888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 34.544 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 141.260000 0.000000 141.640000 0.700000 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7445 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 139.880000 0.000000 140.260000 0.700000 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.837 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 138.500000 0.000000 138.880000 0.700000 ;
    END
  END SS4BEG[0]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.9852 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.761 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met2  ;
    ANTENNAMAXAREACAR 13.2492 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 57.6346 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.694037 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.6396 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.352 LAYER met3  ;
    ANTENNAGATEAREA 1.7067 LAYER met3  ;
    ANTENNAMAXAREACAR 20.8997 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 97.7023 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.694037 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 88.360000 199.560000 88.740000 200.260000 ;
    END
  END S1END[3]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.0314 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 64.652 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 34.8945 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 155.492 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.390645 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.3999 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.928 LAYER met3  ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 52.6969 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 251.052 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.627985 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAGATEAREA 1.7067 LAYER met4  ;
    ANTENNAMAXAREACAR 52.981 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 252.843 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.674423 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 86.520000 199.560000 86.900000 200.260000 ;
    END
  END S1END[2]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4455 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.0346 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.792 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7067 LAYER met4  ;
    ANTENNAMAXAREACAR 56.9262 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 282.651 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.01961 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 85.140000 199.560000 85.520000 200.260000 ;
    END
  END S1END[1]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7881 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5435 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 8.32114 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.8111 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 9.08259 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 27.9457 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.4046 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 120.432 LAYER met4  ;
    ANTENNAGATEAREA 1.7067 LAYER met4  ;
    ANTENNAMAXAREACAR 56.5248 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 296.199 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 83.760000 199.560000 84.140000 200.260000 ;
    END
  END S1END[0]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.0383 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 79.4605 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0707 LAYER met2  ;
    ANTENNAMAXAREACAR 25.384 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 120.481 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.643648 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 1.0707 LAYER met3  ;
    ANTENNAMAXAREACAR 25.6183 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 122.17 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.681007 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.1508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 150.608 LAYER met4  ;
    ANTENNAGATEAREA 1.8132 LAYER met4  ;
    ANTENNAMAXAREACAR 41.1438 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 205.232 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.681007 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 112.740000 199.560000 113.120000 200.260000 ;
    END
  END S2MID[7]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.2209 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.3735 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 24.1447 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 101.611 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.390645 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.9468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.52 LAYER met3  ;
    ANTENNAGATEAREA 1.6542 LAYER met3  ;
    ANTENNAMAXAREACAR 24.7171 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 104.948 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.390645 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 110.900000 199.560000 111.280000 200.260000 ;
    END
  END S2MID[6]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.4737 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.9815 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 26.1951 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 112.194 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.390645 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.8788 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.824 LAYER met3  ;
    ANTENNAGATEAREA 1.8132 LAYER met3  ;
    ANTENNAMAXAREACAR 27.7828 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 120.921 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.390645 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 109.520000 199.560000 109.900000 200.260000 ;
    END
  END S2MID[5]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9755 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.5985 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 13.8077 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 50.2668 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 14.4264 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 54.4813 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.1293 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 274.096 LAYER met4  ;
    ANTENNAGATEAREA 1.6542 LAYER met4  ;
    ANTENNAMAXAREACAR 55.8953 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 287.15 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 108.140000 199.560000 108.520000 200.260000 ;
    END
  END S2MID[4]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7859 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6605 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 11.3573 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.2862 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 13.2298 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 49.3467 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.3938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 279.904 LAYER met4  ;
    ANTENNAGATEAREA 1.8132 LAYER met4  ;
    ANTENNAMAXAREACAR 42.1256 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 203.717 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.381305 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 106.300000 199.560000 106.680000 200.260000 ;
    END
  END S2MID[3]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9297 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3695 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 10.666 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.5583 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.955 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.56 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 26.6655 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 120.963 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.1464 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 162.192 LAYER met4  ;
    ANTENNAGATEAREA 1.6542 LAYER met4  ;
    ANTENNAMAXAREACAR 56.4354 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 284.109 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.80021 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 104.920000 199.560000 105.300000 200.260000 ;
    END
  END S2MID[2]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5499 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.4705 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 11.199 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.2234 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 11.7762 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 41.3826 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.8428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 255.632 LAYER met4  ;
    ANTENNAGATEAREA 1.8132 LAYER met4  ;
    ANTENNAMAXAREACAR 39.3691 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 200.736 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.441028 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 103.540000 199.560000 103.920000 200.260000 ;
    END
  END S2MID[1]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.514 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.301 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 9.46837 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 28.8417 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 10.706 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 36.516 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.3938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 279.904 LAYER met4  ;
    ANTENNAGATEAREA 1.6542 LAYER met4  ;
    ANTENNAMAXAREACAR 45.0271 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 229.167 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.388871 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 101.700000 199.560000 102.080000 200.260000 ;
    END
  END S2MID[0]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8503 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.9825 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 10.6499 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.9045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.127 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.144 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 24.7447 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 111.15 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 45.9937 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 227.656 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.632495 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 100.320000 199.560000 100.700000 200.260000 ;
    END
  END S2END[7]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.0012 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.619 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 26.0353 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 111.62 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.390645 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 26.4883 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 114.706 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.458019 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.4804 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 30.64 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 30.945 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 139.623 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 98.940000 199.560000 99.320000 200.260000 ;
    END
  END S2END[6]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3639 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.6585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1664 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.664 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 7.36531 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 20.6211 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.0676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.968 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 58.8101 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 295.944 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.09371 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 97.560000 199.560000 97.940000 200.260000 ;
    END
  END S2END[5]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6255 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8485 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 10.9333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.8949 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.967 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.624 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 47.6644 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 232.867 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.0686 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 198.64 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 77.8088 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 394.403 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 95.720000 199.560000 96.100000 200.260000 ;
    END
  END S2END[4]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.1947 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.1145 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met2  ;
    ANTENNAMAXAREACAR 21.9836 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 96.2444 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.517922 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 22.79 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 101.165 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.571064 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.4868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.4 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 34.3588 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 168.081 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.571064 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 94.340000 199.560000 94.720000 200.260000 ;
    END
  END S2END[3]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5693 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5775 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 9.44744 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 28.7371 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 10.034 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 32.8963 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.2826 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.448 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 47.2027 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 234.719 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.690147 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 92.960000 199.560000 93.340000 200.260000 ;
    END
  END S2END[2]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5855 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 9.06004 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.6839 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 9.64665 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 30.8431 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.3036 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 258.56 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 75.3428 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 386.438 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 91.120000 199.560000 91.500000 200.260000 ;
    END
  END S2END[1]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1707 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.746 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.3913 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 190.16 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 51.7767 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 265.218 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.910273 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 89.740000 199.560000 90.120000 200.260000 ;
    END
  END S2END[0]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0745 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.9855 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 10.9059 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.758 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 12.1435 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 43.4323 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.2978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 279.392 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 56.5691 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 280.768 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 136.660000 199.560000 137.040000 200.260000 ;
    END
  END S4END[15]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.8557 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.9995 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 16.207 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 62.2636 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.517 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.224 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 31.199 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 143.294 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.2198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 246.976 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 70.4615 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 353.094 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 135.280000 199.560000 135.660000 200.260000 ;
    END
  END S4END[14]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.5613 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.4195 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 12.5484 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.9706 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 13.1671 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 48.185 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.6618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 260 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 54.504 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 269.048 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 133.900000 199.560000 134.280000 200.260000 ;
    END
  END S4END[13]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.3367 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.2865 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 18.6701 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 74.7113 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.54 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.68 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 29.1141 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 131.486 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.5988 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 243.664 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 67.8491 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 338.472 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 132.060000 199.560000 132.440000 200.260000 ;
    END
  END S4END[12]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9833 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.6475 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 17.5118 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 69.0591 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.953 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.216 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 24.305 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 106.363 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.7708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 255.248 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 64.8851 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 323.189 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 130.680000 199.560000 131.060000 200.260000 ;
    END
  END S4END[11]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.1901 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.5535 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 17.4207 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 68.0607 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 18.4997 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 74.8884 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.8188 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 255.504 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 59.1204 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 291.932 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 129.300000 199.560000 129.680000 200.260000 ;
    END
  END S4END[10]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.861 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 11.6133 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.5664 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.111 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.392 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 14.1691 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 54.2708 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.0888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 272.944 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 57.5677 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 286.129 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 127.460000 199.560000 127.840000 200.260000 ;
    END
  END S4END[9]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.2635 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 11.6503 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.7516 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 14.634 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 56.738 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.9298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 256.096 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 55.3491 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 274.285 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 126.080000 199.560000 126.460000 200.260000 ;
    END
  END S4END[8]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.5406 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 127.477 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 32.0662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 142.009 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.170002 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 124.700000 199.560000 125.080000 200.260000 ;
    END
  END S4END[7]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4405 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9335 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 11.2252 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.6259 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 14.0501 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 53.7658 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.3698 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 279.776 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 58.5369 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 291.428 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 123.320000 199.560000 123.700000 200.260000 ;
    END
  END S4END[6]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.9583 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.5125 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 14.4438 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 53.4472 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 15.0625 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 57.6616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.1398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 129.216 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 40.3251 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 208.665 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 121.480000 199.560000 121.860000 200.260000 ;
    END
  END S4END[5]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2563 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.0125 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 11.5839 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.5744 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 13.4564 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 50.6349 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.3068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 263.44 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 55.3412 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 274.42 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 120.100000 199.560000 120.480000 200.260000 ;
    END
  END S4END[4]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.7845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 15.7888 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 60.444 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 17.6614 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 71.5045 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.8048 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 42.096 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 37.0159 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 179.883 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.565409 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 118.720000 199.560000 119.100000 200.260000 ;
    END
  END S4END[3]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.4237 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.7315 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 14.2694 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 52.7306 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 15.6657 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 61.2514 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.6168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 147.76 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 59.8656 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 305.837 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.682809 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 116.880000 199.560000 117.260000 200.260000 ;
    END
  END S4END[2]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6525 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9835 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 10.0283 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.3699 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 11.5834 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 40.7373 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.9426 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 149.968 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 66.459 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 338.883 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 115.500000 199.560000 115.880000 200.260000 ;
    END
  END S4END[1]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6525 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9835 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 11.3616 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.0366 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 11.9482 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 42.1958 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.0096 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 240.992 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 81.5205 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 412.592 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 114.120000 199.560000 114.500000 200.260000 ;
    END
  END S4END[0]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3307 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2665 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 9.56936 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.0752 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.205 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.56 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 16.9423 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 69.4709 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.1258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 267.808 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 59.5228 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 296.967 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 161.040000 199.560000 161.420000 200.260000 ;
    END
  END SS4END[15]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.9834 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 124.691 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 26.5558 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 114.457 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.170002 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 159.660000 199.560000 160.040000 200.260000 ;
    END
  END SS4END[14]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.0253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.7395 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 18.2167 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 72.3119 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.056 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 25.8035 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 113.849 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.2198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 230.976 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 62.5176 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 310.057 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 157.820000 199.560000 158.200000 200.260000 ;
    END
  END SS4END[13]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.5663 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.4445 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 23.7992 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 100.38 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 27.1003 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 119.059 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.9128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 202.672 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 59.3062 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 291.224 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 156.440000 199.560000 156.820000 200.260000 ;
    END
  END SS4END[12]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.7848 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.655 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 15.4329 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 58.6646 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.61 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.72 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 30.6388 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 140.836 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.2828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 247.312 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 69.9548 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 350.921 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 155.060000 199.560000 155.440000 200.260000 ;
    END
  END SS4END[11]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8487 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.8565 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 10.761 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.0334 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.592 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.624 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 12.1228 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 43.3701 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.3438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 258.304 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 53.1896 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 262.793 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 153.680000 199.560000 154.060000 200.260000 ;
    END
  END SS4END[10]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5621 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4235 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 8.54198 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.9383 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 10.2558 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 34.1523 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.9798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 261.696 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 51.8628 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 267.715 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 151.840000 199.560000 152.220000 200.260000 ;
    END
  END SS4END[9]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.8809 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.1255 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 33.8496 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 150.476 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.584 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 40.8015 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 188.627 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.2288 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 183.024 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 69.8779 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 344.101 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.460000 199.560000 150.840000 200.260000 ;
    END
  END SS4END[8]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.9066 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 139.307 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 30.783 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 135.593 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.170002 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 149.080000 199.560000 149.460000 200.260000 ;
    END
  END SS4END[7]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.8941 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.0835 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 15.3515 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 58.1412 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 15.9381 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 62.3004 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.0478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 219.392 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 50.8071 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 248.668 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 147.240000 199.560000 147.620000 200.260000 ;
    END
  END SS4END[6]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6411 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2279 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.992 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 9.52818 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 31.3274 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.9668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 282.96 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 54.5221 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 271.694 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 145.860000 199.560000 146.240000 200.260000 ;
    END
  END SS4END[5]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4139 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.6725 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 12.905 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 45.6372 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 15.4125 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 60.084 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.1128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 273.072 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 58.8314 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 292.051 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 144.480000 199.560000 144.860000 200.260000 ;
    END
  END SS4END[4]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.0116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 79.016 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met2  ;
    ANTENNAMAXAREACAR 22.8297 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 105.247 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.46478 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 142.640000 199.560000 143.020000 200.260000 ;
    END
  END SS4END[3]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1316 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.379 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 19.3181 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.8192 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.091 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.952 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 26.4288 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 116.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 100.912 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 82.2555 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 412.196 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.632495 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 141.260000 199.560000 141.640000 200.260000 ;
    END
  END SS4END[2]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.971 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.059 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met2  ;
    ANTENNAMAXAREACAR 33.2867 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 147.851 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 139.880000 199.560000 140.260000 200.260000 ;
    END
  END SS4END[1]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7148 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.016 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 15.3501 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 57.5857 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.655 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.408 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 16.8569 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 67.726 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.486312 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.8876 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 235.008 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 83.6263 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 430.466 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 138.500000 199.560000 138.880000 200.260000 ;
    END
  END SS4END[0]
  PIN W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 9.350000 0.700000 9.730000 ;
    END
  END W1BEG[3]
  PIN W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.36 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 7.520000 0.700000 7.900000 ;
    END
  END W1BEG[2]
  PIN W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 6.300000 0.700000 6.680000 ;
    END
  END W1BEG[1]
  PIN W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 5.080000 0.700000 5.460000 ;
    END
  END W1BEG[0]
  PIN W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 20.940000 0.700000 21.320000 ;
    END
  END W2BEG[7]
  PIN W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.712 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 19.720000 0.700000 20.100000 ;
    END
  END W2BEG[6]
  PIN W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 17.890000 0.700000 18.270000 ;
    END
  END W2BEG[5]
  PIN W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.2644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.072 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 16.670000 0.700000 17.050000 ;
    END
  END W2BEG[4]
  PIN W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 15.450000 0.700000 15.830000 ;
    END
  END W2BEG[3]
  PIN W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.677 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 13.620000 0.700000 14.000000 ;
    END
  END W2BEG[2]
  PIN W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.1304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.024 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 12.400000 0.700000 12.780000 ;
    END
  END W2BEG[1]
  PIN W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 10.570000 0.700000 10.950000 ;
    END
  END W2BEG[0]
  PIN W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 33.140000 0.700000 33.520000 ;
    END
  END W2BEGb[7]
  PIN W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 31.310000 0.700000 31.690000 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.4426 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 30.090000 0.700000 30.470000 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 28.870000 0.700000 29.250000 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 27.040000 0.700000 27.420000 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 37.7776 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 201.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 25.820000 0.700000 26.200000 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 23.990000 0.700000 24.370000 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 22.770000 0.700000 23.150000 ;
    END
  END W2BEGb[0]
  PIN WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.8638 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.744 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 56.930000 0.700000 57.310000 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 55.100000 0.700000 55.480000 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 53.880000 0.700000 54.260000 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.5224 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.448 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 52.660000 0.700000 53.040000 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2654 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.744 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 50.830000 0.700000 51.210000 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.1964 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.376 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 49.610000 0.700000 49.990000 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 47.780000 0.700000 48.160000 ;
    END
  END WW4BEG[9]
  PIN WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.656 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 46.560000 0.700000 46.940000 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 44.730000 0.700000 45.110000 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 43.510000 0.700000 43.890000 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.4024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.808 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 42.290000 0.700000 42.670000 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 40.460000 0.700000 40.840000 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.0584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 39.240000 0.700000 39.620000 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 37.410000 0.700000 37.790000 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 36.190000 0.700000 36.570000 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 34.360000 0.700000 34.740000 ;
    END
  END WW4BEG[0]
  PIN W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 74.620000 0.700000 75.000000 ;
    END
  END W6BEG[11]
  PIN W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 73.400000 0.700000 73.780000 ;
    END
  END W6BEG[10]
  PIN W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 71.570000 0.700000 71.950000 ;
    END
  END W6BEG[9]
  PIN W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 70.350000 0.700000 70.730000 ;
    END
  END W6BEG[8]
  PIN W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.5404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.544 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 68.520000 0.700000 68.900000 ;
    END
  END W6BEG[7]
  PIN W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 67.300000 0.700000 67.680000 ;
    END
  END W6BEG[6]
  PIN W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.3684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.96 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 66.080000 0.700000 66.460000 ;
    END
  END W6BEG[5]
  PIN W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 64.250000 0.700000 64.630000 ;
    END
  END W6BEG[4]
  PIN W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 63.030000 0.700000 63.410000 ;
    END
  END W6BEG[3]
  PIN W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 61.200000 0.700000 61.580000 ;
    END
  END W6BEG[2]
  PIN W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 59.980000 0.700000 60.360000 ;
    END
  END W6BEG[1]
  PIN W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 58.150000 0.700000 58.530000 ;
    END
  END W6BEG[0]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.9752 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 144.8 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 58.3612 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 299.935 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.893789 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 65.9973 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 355.744 LAYER met4  ;
    ANTENNAGATEAREA 2.1837 LAYER met4  ;
    ANTENNAMAXAREACAR 88.5839 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 462.844 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 9.350000 200.100000 9.730000 ;
    END
  END W1END[3]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.9304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.424 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 74.5632 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 367.088 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.666902 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.5838 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 195.584 LAYER met4  ;
    ANTENNAGATEAREA 2.1837 LAYER met4  ;
    ANTENNAMAXAREACAR 91.3163 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 456.653 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.851572 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 7.520000 200.100000 7.900000 ;
    END
  END W1END[2]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.1474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.248 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 24.8753 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 119.595 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.666902 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.3294 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 131.168 LAYER met4  ;
    ANTENNAGATEAREA 1.8657 LAYER met4  ;
    ANTENNAMAXAREACAR 65.9112 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 333.322 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.742558 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 6.300000 200.100000 6.680000 ;
    END
  END W1END[1]
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.781 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.632 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 21.7295 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 93.7037 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.6316 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 62.976 LAYER met4  ;
    ANTENNAGATEAREA 1.7067 LAYER met4  ;
    ANTENNAMAXAREACAR 41.3342 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 202.389 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.527673 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 5.080000 200.100000 5.460000 ;
    END
  END W1END[0]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7526 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.3515 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 104.144 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8132 LAYER met4  ;
    ANTENNAMAXAREACAR 64.0066 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 340.89 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 20.940000 200.100000 21.320000 ;
    END
  END W2MID[7]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 27.0874 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 144.928 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 70.2563 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 354.47 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.1522 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 300.88 LAYER met4  ;
    ANTENNAGATEAREA 1.6542 LAYER met4  ;
    ANTENNAMAXAREACAR 104.201 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 536.358 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 19.720000 200.100000 20.100000 ;
    END
  END W2MID[6]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.8818 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.84 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8132 LAYER met3  ;
    ANTENNAMAXAREACAR 24.5444 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 120.665 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 17.890000 200.100000 18.270000 ;
    END
  END W2MID[5]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 34.3482 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 183.656 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6542 LAYER met3  ;
    ANTENNAMAXAREACAR 40.9732 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 205.009 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.49758 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 16.670000 200.100000 17.050000 ;
    END
  END W2MID[4]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 51.5952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 275.64 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8132 LAYER met3  ;
    ANTENNAMAXAREACAR 38.7965 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 197.913 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.493797 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 15.450000 200.100000 15.830000 ;
    END
  END W2MID[3]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.6649 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.008 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 20.7898 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 87.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.388016 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.2948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 71.376 LAYER met4  ;
    ANTENNAGATEAREA 1.6542 LAYER met4  ;
    ANTENNAMAXAREACAR 51.2367 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 256.533 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.632495 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 13.620000 200.100000 14.000000 ;
    END
  END W2MID[2]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.105 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.36 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 34.6151 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 163.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.5524 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.024 LAYER met4  ;
    ANTENNAGATEAREA 1.8132 LAYER met4  ;
    ANTENNAMAXAREACAR 44.8252 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 229.979 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.0123 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 12.400000 200.100000 12.780000 ;
    END
  END W2MID[1]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 33.87 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 181.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6542 LAYER met3  ;
    ANTENNAMAXAREACAR 36.0101 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 178.846 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.632495 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 10.570000 200.100000 10.950000 ;
    END
  END W2MID[0]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.6324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.168 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 37.4375 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 175.342 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.5108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.528 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 47.4841 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 242.229 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.490985 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 33.140000 200.100000 33.520000 ;
    END
  END W2END[7]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.8882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 138.536 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 65.6754 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 321.815 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 31.310000 200.100000 31.690000 ;
    END
  END W2END[6]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 15.0752 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 57.8836 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.3026 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 55.888 LAYER met4  ;
    ANTENNAGATEAREA 0.7527 LAYER met4  ;
    ANTENNAMAXAREACAR 33.9855 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 171.28 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 30.090000 200.100000 30.470000 ;
    END
  END W2END[5]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 34.231 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 183.032 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 93.4755 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 475.845 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.6938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.504 LAYER met4  ;
    ANTENNAGATEAREA 1.5477 LAYER met4  ;
    ANTENNAMAXAREACAR 96.5083 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 492.324 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.678167 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 28.870000 200.100000 29.250000 ;
    END
  END W2END[4]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.7614 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 121.856 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 80.2011 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 400.605 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.4466 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.656 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 83.403 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 418.36 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.942767 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 27.040000 200.100000 27.420000 ;
    END
  END W2END[3]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 29.9614 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 160.256 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 82.3734 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 417.259 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.0216 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 49.056 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 88.8698 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 452.584 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 25.820000 200.100000 26.200000 ;
    END
  END W2END[2]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 29.7378 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 159.072 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met3  ;
    ANTENNAMAXAREACAR 41.9567 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 211.223 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.506709 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 23.990000 200.100000 24.370000 ;
    END
  END W2END[1]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.9804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 139.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 71.8627 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 361.452 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.512537 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    ANTENNAGATEAREA 0.7527 LAYER met4  ;
    ANTENNAMAXAREACAR 72.993 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 368.105 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 22.770000 200.100000 23.150000 ;
    END
  END W2END[0]
  PIN WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 53.6598 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 286.656 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 54.7719 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 270.682 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 56.930000 200.100000 57.310000 ;
    END
  END WW4END[15]
  PIN WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.8653 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.072 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 47.7709 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 236.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.343 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 78.848 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 59.9549 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 303.46 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 55.100000 200.100000 55.480000 ;
    END
  END WW4END[14]
  PIN WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 53.2542 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 284.488 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 54.6077 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 269.597 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 53.880000 200.100000 54.260000 ;
    END
  END WW4END[13]
  PIN WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 36.7234 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 196.32 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 93.6759 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 478.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.888 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 95.1759 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 486.81 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 52.660000 200.100000 53.040000 ;
    END
  END WW4END[12]
  PIN WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 51.0798 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 272.896 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 54.9166 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 270.571 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 50.830000 200.100000 51.210000 ;
    END
  END WW4END[11]
  PIN WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 54.3582 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 290.376 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 55.3297 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 273.52 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 49.610000 200.100000 49.990000 ;
    END
  END WW4END[10]
  PIN WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.39 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.88 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 27.1946 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 123.329 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 62.0398 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 329.993 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 47.780000 200.100000 48.160000 ;
    END
  END WW4END[9]
  PIN WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 52.1952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 278.84 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 55.4914 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 273.736 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 46.560000 200.100000 46.940000 ;
    END
  END WW4END[8]
  PIN WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 49.6504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 265.264 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 121.205 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 626.513 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 122.083 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 631.596 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 44.730000 200.100000 45.110000 ;
    END
  END WW4END[7]
  PIN WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 46.7262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 249.672 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 57.3425 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 281.423 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 43.510000 200.100000 43.890000 ;
    END
  END WW4END[6]
  PIN WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.4045 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.144 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 13.553 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 52.0704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.6654 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 68.96 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 49.2226 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 262.413 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 42.290000 200.100000 42.670000 ;
    END
  END WW4END[5]
  PIN WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 50.7108 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 270.928 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 57.5003 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 283.344 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 40.460000 200.100000 40.840000 ;
    END
  END WW4END[4]
  PIN WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.8462 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 56.3528 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 284.563 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.407128 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 39.240000 200.100000 39.620000 ;
    END
  END WW4END[3]
  PIN WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7736 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.6937 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 129.184 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0707 LAYER met4  ;
    ANTENNAMAXAREACAR 69.2883 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 354.625 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 37.410000 200.100000 37.790000 ;
    END
  END WW4END[2]
  PIN WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 31.6153 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 169.072 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 63.0569 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 315.044 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.642217 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.3948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.576 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 86.5238 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 440.717 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.642217 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 36.190000 200.100000 36.570000 ;
    END
  END WW4END[1]
  PIN WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.1938 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 61.8734 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 308.257 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.548637 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 34.360000 200.100000 34.740000 ;
    END
  END WW4END[0]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.4013 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.264 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 51.8995 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 257.918 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 52.4667 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 261.343 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 74.620000 200.100000 75.000000 ;
    END
  END W6END[11]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 24.064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 128.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 72.7518 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 364.617 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.1578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.312 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 77.9827 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 392.915 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 73.400000 200.100000 73.780000 ;
    END
  END W6END[10]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 55.9692 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 298.968 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 52.8689 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 262.099 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 71.570000 200.100000 71.950000 ;
    END
  END W6END[9]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 53.5564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 286.096 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 135.616 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 701.295 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 136.339 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 705.549 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 70.350000 200.100000 70.730000 ;
    END
  END W6END[8]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.1785 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.272 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 21.6273 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 95.4911 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 68.3288 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 363.658 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 68.520000 200.100000 68.900000 ;
    END
  END W6END[7]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 10.6243 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 35.7442 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.3486 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.8 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 36.6283 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 195.029 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 67.300000 200.100000 67.680000 ;
    END
  END W6END[6]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 39.9715 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 213.168 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 97.219 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 498.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.8256 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.344 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 103.017 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 530.163 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 66.080000 200.100000 66.460000 ;
    END
  END W6END[5]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 50.2662 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 268.552 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 57.4182 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 282.524 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.42052 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 64.250000 200.100000 64.630000 ;
    END
  END W6END[4]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 53.7102 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 286.92 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 52.6141 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 259.779 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 63.030000 200.100000 63.410000 ;
    END
  END W6END[3]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5874 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 66.6499 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 230.798 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.512537 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.5966 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 89.456 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 80.7482 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 306.789 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.512537 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 61.200000 200.100000 61.580000 ;
    END
  END W6END[2]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.9634 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 27.425 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 122.726 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.525393 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.6097 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 78.384 LAYER met4  ;
    ANTENNAGATEAREA 2.0247 LAYER met4  ;
    ANTENNAMAXAREACAR 34.6407 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 165.517 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.779245 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 59.980000 200.100000 60.360000 ;
    END
  END W6END[1]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 27.166 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 146.288 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met3  ;
    ANTENNAMAXAREACAR 50.1129 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 251.156 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.665023 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.936 LAYER met4  ;
    ANTENNAGATEAREA 1.7067 LAYER met4  ;
    ANTENNAMAXAREACAR 50.9331 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 255.806 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.665023 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 58.150000 200.100000 58.530000 ;
    END
  END W6END[0]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.2515 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.1947 LAYER met3  ;
    ANTENNAMAXAREACAR 23.6109 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 116.613 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 162.420000 0.000000 162.800000 0.700000 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1275 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.6275 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 162.420000 199.560000 162.800000 200.260000 ;
    END
  END UserCLKo
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.6814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.744 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 31.4143 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 145.963 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.7614 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 244.992 LAYER met4  ;
    ANTENNAGATEAREA 3.4932 LAYER met4  ;
    ANTENNAMAXAREACAR 60.0605 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 309.536 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.00269 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 194.180000 0.700000 194.560000 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.94 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.48 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 22.1148 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 109.169 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.525393 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.2178 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 275.504 LAYER met4  ;
    ANTENNAGATEAREA 3.4932 LAYER met4  ;
    ANTENNAMAXAREACAR 60.1602 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 307.737 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 192.350000 0.700000 192.730000 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.153 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 139.936 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 68.9312 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 347.108 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.486312 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.9956 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 285.936 LAYER met4  ;
    ANTENNAGATEAREA 3.3342 LAYER met4  ;
    ANTENNAMAXAREACAR 84.8258 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 432.867 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.884067 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 191.130000 0.700000 191.510000 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.2854 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.984 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 16.0939 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 65.5349 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.5194 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 94.848 LAYER met4  ;
    ANTENNAGATEAREA 3.4932 LAYER met4  ;
    ANTENNAMAXAREACAR 62.4446 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 311.687 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.87673 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 189.300000 0.700000 189.680000 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.1926 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.8766 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 85.136 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4932 LAYER met4  ;
    ANTENNAMAXAREACAR 58.8782 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 297.791 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.6587 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 188.080000 0.700000 188.460000 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.9285 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 90.272 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 44.1049 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 215.355 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.4126 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 303.68 LAYER met4  ;
    ANTENNAGATEAREA 3.4932 LAYER met4  ;
    ANTENNAMAXAREACAR 60.2542 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 302.29 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 186.250000 0.700000 186.630000 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.5964 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.976 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 28.4307 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 142.721 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.624206 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 64.5837 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 349.136 LAYER met4  ;
    ANTENNAGATEAREA 3.6522 LAYER met4  ;
    ANTENNAMAXAREACAR 56.9741 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 294.258 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.854717 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 185.030000 0.700000 185.410000 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8237 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.272 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 12.8698 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 49.3186 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.542641 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.7199 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 267.52 LAYER met4  ;
    ANTENNAGATEAREA 3.8112 LAYER met4  ;
    ANTENNAMAXAREACAR 76.4329 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 394.752 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.99413 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 183.200000 0.700000 183.580000 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.9367 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.384 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 22.2324 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 94.753 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.05567 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.5692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 303.584 LAYER met4  ;
    ANTENNAGATEAREA 3.8112 LAYER met4  ;
    ANTENNAMAXAREACAR 72.087 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 361.224 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.09371 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 181.980000 0.700000 182.360000 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.926 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1752 LAYER met3  ;
    ANTENNAMAXAREACAR 41.2132 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 202.119 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.830015 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.3656 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 104.224 LAYER met4  ;
    ANTENNAGATEAREA 3.8112 LAYER met4  ;
    ANTENNAMAXAREACAR 46.2945 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 229.466 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.830015 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 180.760000 0.700000 181.140000 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 43.2023 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 231.336 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 57.4378 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 290.161 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.585325 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 66.1728 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 354.784 LAYER met4  ;
    ANTENNAGATEAREA 3.8112 LAYER met4  ;
    ANTENNAMAXAREACAR 74.8006 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 383.251 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.938933 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 178.930000 0.700000 179.310000 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.536 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 70.8346 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 369.497 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.2195 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.4023 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 277.424 LAYER met4  ;
    ANTENNAGATEAREA 3.8112 LAYER met4  ;
    ANTENNAMAXAREACAR 91.957 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 483.631 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.2195 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 177.710000 0.700000 178.090000 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 20.7702 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 100.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.666902 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.3425 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 136.096 LAYER met4  ;
    ANTENNAGATEAREA 3.8112 LAYER met4  ;
    ANTENNAMAXAREACAR 65.2521 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 331.303 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.862354 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 175.880000 0.700000 176.260000 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.3966 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.5249 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 282 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8112 LAYER met4  ;
    ANTENNAMAXAREACAR 65.0151 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 344.452 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 174.660000 0.700000 175.040000 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8216 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.04 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.3007 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 206.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8112 LAYER met4  ;
    ANTENNAMAXAREACAR 68.1082 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 361.676 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 172.830000 0.700000 173.210000 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.3694 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.432 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 39.3455 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 198.244 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.642217 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.3909 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 260.432 LAYER met4  ;
    ANTENNAGATEAREA 3.8112 LAYER met4  ;
    ANTENNAMAXAREACAR 89.1587 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 472.761 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 171.610000 0.700000 171.990000 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.8714 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.776 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6982 LAYER met3  ;
    ANTENNAMAXAREACAR 34.8453 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 169.75 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.509254 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.3274 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 109.824 LAYER met4  ;
    ANTENNAGATEAREA 3.8112 LAYER met4  ;
    ANTENNAMAXAREACAR 52.8035 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 266.037 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 169.780000 0.700000 170.160000 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 23.4866 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 127.12 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7067 LAYER met3  ;
    ANTENNAMAXAREACAR 38.1765 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 190.973 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.655932 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.2991 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 147.472 LAYER met4  ;
    ANTENNAGATEAREA 3.8112 LAYER met4  ;
    ANTENNAMAXAREACAR 62.7042 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 322.193 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.0398 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 168.560000 0.700000 168.940000 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.6561 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.928 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met3  ;
    ANTENNAMAXAREACAR 51.4524 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 256.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.665023 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.3242 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 120.944 LAYER met4  ;
    ANTENNAGATEAREA 3.8112 LAYER met4  ;
    ANTENNAMAXAREACAR 84.3731 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 439.943 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.12342 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 167.340000 0.700000 167.720000 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.9793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.68 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0707 LAYER met3  ;
    ANTENNAMAXAREACAR 28.1073 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 136.585 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.585996 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.7753 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 96.208 LAYER met4  ;
    ANTENNAGATEAREA 3.8112 LAYER met4  ;
    ANTENNAMAXAREACAR 50.7851 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 257.307 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.646721 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 165.510000 0.700000 165.890000 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.0049 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.664 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 25.0076 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 118.842 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.642217 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.4942 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 111.184 LAYER met4  ;
    ANTENNAGATEAREA 3.8112 LAYER met4  ;
    ANTENNAMAXAREACAR 84.9794 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 440.747 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.871843 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 164.290000 0.700000 164.670000 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.4952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 40.2824 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 199.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.769494 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 64.641 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 346.624 LAYER met4  ;
    ANTENNAGATEAREA 3.8112 LAYER met4  ;
    ANTENNAMAXAREACAR 89.2052 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 462.425 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.13564 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 162.460000 0.700000 162.840000 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 134.912 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5477 LAYER met3  ;
    ANTENNAMAXAREACAR 54.1542 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 271.972 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.878105 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 97.6533 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 524.096 LAYER met4  ;
    ANTENNAGATEAREA 3.8112 LAYER met4  ;
    ANTENNAMAXAREACAR 90.9202 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 479.04 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 161.240000 0.700000 161.620000 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.4942 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 116.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5477 LAYER met3  ;
    ANTENNAMAXAREACAR 44.1117 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 220.118 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.993769 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.8058 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 119.12 LAYER met4  ;
    ANTENNAGATEAREA 3.8112 LAYER met4  ;
    ANTENNAMAXAREACAR 72.3272 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 378.318 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.72264 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 159.410000 0.700000 159.790000 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.4681 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.432 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met3  ;
    ANTENNAMAXAREACAR 29.4262 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 145.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.661299 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.6489 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 117.808 LAYER met4  ;
    ANTENNAGATEAREA 3.8112 LAYER met4  ;
    ANTENNAMAXAREACAR 56.478 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 282.573 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.01824 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 158.190000 0.700000 158.570000 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.2222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.784 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0707 LAYER met3  ;
    ANTENNAMAXAREACAR 31.1236 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 155.102 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.612202 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 58.8279 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 318.448 LAYER met4  ;
    ANTENNAGATEAREA 3.6522 LAYER met4  ;
    ANTENNAMAXAREACAR 90.9836 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 482.269 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.58113 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 156.360000 0.700000 156.740000 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.9306 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.088 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 32.0004 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 148.842 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.527053 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.2475 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 228.608 LAYER met4  ;
    ANTENNAGATEAREA 3.8112 LAYER met4  ;
    ANTENNAMAXAREACAR 65.4313 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 334.485 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 155.140000 0.700000 155.520000 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 14.6299 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 56.6103 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.512537 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.3137 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 265.824 LAYER met4  ;
    ANTENNAGATEAREA 3.8112 LAYER met4  ;
    ANTENNAMAXAREACAR 75.1743 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 398.252 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.2195 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 153.920000 0.700000 154.300000 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.66358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.128 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 47.229 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 236.286 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.0353 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.361 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 174.464 LAYER met4  ;
    ANTENNAGATEAREA 3.6522 LAYER met4  ;
    ANTENNAMAXAREACAR 56.0897 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 284.055 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.0353 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 152.090000 0.700000 152.470000 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4766 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 54.3252 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 291.616 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4932 LAYER met4  ;
    ANTENNAMAXAREACAR 68.3263 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 345.765 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.660197 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 150.870000 0.700000 151.250000 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9276 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.3805 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 223.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4932 LAYER met4  ;
    ANTENNAMAXAREACAR 52.9413 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 269.548 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 149.040000 0.700000 149.420000 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.008 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 18.771 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 78.1633 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.459679 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.6548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.296 LAYER met4  ;
    ANTENNAGATEAREA 3.1752 LAYER met4  ;
    ANTENNAMAXAREACAR 62.5883 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 310.628 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.731847 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 147.820000 0.700000 148.200000 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.4364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.656 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 194.180000 200.100000 194.560000 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 192.350000 200.100000 192.730000 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.8614 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.256 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 191.130000 200.100000 191.510000 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 189.300000 200.100000 189.680000 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.3704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.304 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 188.080000 200.100000 188.460000 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 186.250000 200.100000 186.630000 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 185.030000 200.100000 185.410000 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 183.200000 200.100000 183.580000 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.0598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.456 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 181.980000 200.100000 182.360000 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 180.760000 200.100000 181.140000 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 178.930000 200.100000 179.310000 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.8734 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.32 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 177.710000 200.100000 178.090000 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 175.880000 200.100000 176.260000 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 174.660000 200.100000 175.040000 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 172.830000 200.100000 173.210000 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.7484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.32 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 171.610000 200.100000 171.990000 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 169.780000 200.100000 170.160000 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 168.560000 200.100000 168.940000 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.4944 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.632 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 167.340000 200.100000 167.720000 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4634 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 165.510000 200.100000 165.890000 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.3684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.96 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 164.290000 200.100000 164.670000 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.9294 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.952 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 162.460000 200.100000 162.840000 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 161.240000 200.100000 161.620000 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8334 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.152 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 159.410000 200.100000 159.790000 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 158.190000 200.100000 158.570000 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.6784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 156.360000 200.100000 156.740000 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 155.140000 200.100000 155.520000 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.3754 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.096 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 153.920000 200.100000 154.300000 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 152.090000 200.100000 152.470000 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7574 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.368 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 150.870000 200.100000 151.250000 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.2644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.072 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 149.040000 200.100000 149.420000 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.5404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.544 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 147.820000 200.100000 148.200000 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.5228 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.066 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 12.1969 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.9979 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 116.816 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 62.1808 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 310.726 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.486312 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.6884 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 234.416 LAYER met4  ;
    ANTENNAGATEAREA 4.4472 LAYER met4  ;
    ANTENNAMAXAREACAR 72.0046 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 363.437 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.745949 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 194.160000 0.000000 194.540000 0.700000 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 29.1398 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 142.751 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.7192 LAYER met2  ;
    ANTENNAMAXAREACAR 21.0649 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 96.0889 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.46478 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 192.780000 0.000000 193.160000 0.700000 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.7491 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.7985 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met2  ;
    ANTENNAMAXAREACAR 22.9148 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 104.405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.497308 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.0115 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.664 LAYER met3  ;
    ANTENNAGATEAREA 5.7192 LAYER met3  ;
    ANTENNAMAXAREACAR 30.0401 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 144.537 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.625641 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 191.400000 0.000000 191.780000 0.700000 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.2508 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 74.9 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7067 LAYER met2  ;
    ANTENNAMAXAREACAR 25.8541 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 122.814 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.653163 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3871 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.608 LAYER met3  ;
    ANTENNAGATEAREA 5.7192 LAYER met3  ;
    ANTENNAMAXAREACAR 27.8451 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 133.761 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.653459 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 190.020000 0.000000 190.400000 0.700000 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.0304 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.549 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met2  ;
    ANTENNAMAXAREACAR 12.4803 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.6105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.367145 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.3575 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.176 LAYER met3  ;
    ANTENNAGATEAREA 5.7192 LAYER met3  ;
    ANTENNAMAXAREACAR 29.3462 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 141.131 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.641057 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 188.180000 0.000000 188.560000 0.700000 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.957 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 7.66483 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.824 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.0173 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.632 LAYER met3  ;
    ANTENNAGATEAREA 3.2967 LAYER met3  ;
    ANTENNAMAXAREACAR 26.8838 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 130.219 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.6903 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.1217 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.448 LAYER met4  ;
    ANTENNAGATEAREA 5.7192 LAYER met4  ;
    ANTENNAMAXAREACAR 36.325 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 178.347 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.6903 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 186.800000 0.000000 187.180000 0.700000 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.0916 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 122.542 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1377 LAYER met2  ;
    ANTENNAMAXAREACAR 17.1478 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 79.8566 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.490276 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.25537 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.872 LAYER met3  ;
    ANTENNAGATEAREA 3.1377 LAYER met3  ;
    ANTENNAMAXAREACAR 18.8227 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 89.0583 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.528521 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.1472 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 184 LAYER met4  ;
    ANTENNAGATEAREA 5.7192 LAYER met4  ;
    ANTENNAMAXAREACAR 38.1323 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 188.078 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 185.420000 0.000000 185.800000 0.700000 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0137 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.992 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.7192 LAYER met3  ;
    ANTENNAMAXAREACAR 38.162 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 185.15 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.471774 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 183.580000 0.000000 183.960000 0.700000 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8323 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8535 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 8.7504 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.1622 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 28.291 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 153.704 LAYER met3  ;
    ANTENNAGATEAREA 5.5602 LAYER met3  ;
    ANTENNAMAXAREACAR 29.9469 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 145.851 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.59776 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    ANTENNAGATEAREA 5.7192 LAYER met4  ;
    ANTENNAMAXAREACAR 30.2236 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 147.41 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 182.200000 0.000000 182.580000 0.700000 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.8059 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 83.6325 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 34.3756 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 163.222 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.532154 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.69 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.48 LAYER met3  ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 47.3283 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 233.089 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.599528 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 132.528 LAYER met4  ;
    ANTENNAGATEAREA 5.7192 LAYER met4  ;
    ANTENNAMAXAREACAR 51.596 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 256.261 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.942894 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 180.820000 0.000000 181.200000 0.700000 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.2691 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.4965 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met2  ;
    ANTENNAMAXAREACAR 31.8026 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 139.826 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.376412 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.8878 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.672 LAYER met3  ;
    ANTENNAGATEAREA 5.3637 LAYER met3  ;
    ANTENNAMAXAREACAR 33.0868 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 146.849 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.631097 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.3278 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.552 LAYER met4  ;
    ANTENNAGATEAREA 5.7192 LAYER met4  ;
    ANTENNAMAXAREACAR 35.02 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 181.718 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.68736 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 179.440000 0.000000 179.820000 0.700000 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.6158 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.536 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 18.9354 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 79.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.4872 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 196.48 LAYER met4  ;
    ANTENNAGATEAREA 5.7192 LAYER met4  ;
    ANTENNAMAXAREACAR 57.0628 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 300.612 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 177.600000 0.000000 177.980000 0.700000 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7179 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3105 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 12.4743 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.6002 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 13.5533 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 50.4279 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.4028 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 231.952 LAYER met4  ;
    ANTENNAGATEAREA 5.7192 LAYER met4  ;
    ANTENNAMAXAREACAR 46.3086 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 230.136 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.975494 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 176.220000 0.000000 176.600000 0.700000 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.9289 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 133.913 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9492 LAYER met2  ;
    ANTENNAMAXAREACAR 34.0921 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 165.131 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.506921 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.7786 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.56 LAYER met3  ;
    ANTENNAGATEAREA 5.5602 LAYER met3  ;
    ANTENNAMAXAREACAR 55.1433 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 270.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.582037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.888 LAYER met4  ;
    ANTENNAGATEAREA 5.7192 LAYER met4  ;
    ANTENNAMAXAREACAR 55.452 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 272.289 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 174.840000 0.000000 175.220000 0.700000 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.2551 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.9965 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 14.6821 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 54.6388 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 18.4594 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 75.8581 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 55.1616 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 295.136 LAYER met4  ;
    ANTENNAGATEAREA 5.7192 LAYER met4  ;
    ANTENNAMAXAREACAR 48.1303 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 242.903 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.803144 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 173.000000 0.000000 173.380000 0.700000 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2975 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 7.84173 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.6855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 10.6667 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 36.8254 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 85.3584 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 458.528 LAYER met4  ;
    ANTENNAGATEAREA 5.7192 LAYER met4  ;
    ANTENNAMAXAREACAR 51.7676 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 273.685 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.19033 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 171.620000 0.000000 172.000000 0.700000 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.0527 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.7485 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 36.5123 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 172.295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.532154 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.6082 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.248 LAYER met3  ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 39.2211 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 179.45 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.599528 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.5983 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 191.264 LAYER met4  ;
    ANTENNAGATEAREA 5.5602 LAYER met4  ;
    ANTENNAMAXAREACAR 49.4615 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 241.957 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 170.240000 0.000000 170.620000 0.700000 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2599 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.561 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 12.0032 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.4359 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.706 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.68 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 41.2326 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 198.43 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.486312 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 73.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 398.56 LAYER met4  ;
    ANTENNAGATEAREA 5.0832 LAYER met4  ;
    ANTENNAMAXAREACAR 55.7604 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 276.837 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 168.400000 0.000000 168.780000 0.700000 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.0984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.968 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 14.0083 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 55.1622 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.7251 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 309.744 LAYER met4  ;
    ANTENNAGATEAREA 5.2422 LAYER met4  ;
    ANTENNAMAXAREACAR 47.9003 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 239.975 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.990795 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 167.020000 0.000000 167.400000 0.700000 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3245 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.1685 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 9.5551 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 28.8498 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 10.4753 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 34.8309 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.5712 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 324.928 LAYER met4  ;
    ANTENNAGATEAREA 4.4472 LAYER met4  ;
    ANTENNAMAXAREACAR 52.0425 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 262.988 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.19033 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 165.640000 0.000000 166.020000 0.700000 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4622 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.203 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 194.160000 199.560000 194.540000 200.260000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2982 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.265 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 192.780000 199.560000 193.160000 200.260000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.6038 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.911 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 191.400000 199.560000 191.780000 200.260000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.3994 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.889 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 190.020000 199.560000 190.400000 200.260000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.7022 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.403 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 188.180000 199.560000 188.560000 200.260000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.5458 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.048 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 186.800000 199.560000 187.180000 200.260000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7898 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.723 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 185.420000 199.560000 185.800000 200.260000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6218 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.001 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 183.580000 199.560000 183.960000 200.260000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8114 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.949 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 182.200000 199.560000 182.580000 200.260000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.067 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.227 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 180.820000 199.560000 181.200000 200.260000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3834 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.809 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 179.440000 199.560000 179.820000 200.260000 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.751 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 177.600000 199.560000 177.980000 200.260000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.427 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.909 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 176.220000 199.560000 176.600000 200.260000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.893 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.357 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 174.840000 199.560000 175.220000 200.260000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1766 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.775 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 173.000000 199.560000 173.380000 200.260000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.955 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.667 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 171.620000 199.560000 172.000000 200.260000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2094 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.939 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 170.240000 199.560000 170.620000 200.260000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5574 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.679 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 168.400000 199.560000 168.780000 200.260000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1766 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.775 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 167.020000 199.560000 167.400000 200.260000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5574 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.679 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 165.640000 199.560000 166.020000 200.260000 ;
    END
  END FrameStrobe_O[0]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 198.900000 195.020000 200.100000 196.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 195.020000 1.200000 196.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.900000 2.850000 200.100000 4.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 1.200000 4.050000 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.070000 199.060000 197.270000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.070000 0.000000 197.270000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 199.060000 4.030000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 0.000000 4.030000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 200.100000 4.050000 ;
        RECT 0.000000 195.020000 200.100000 196.220000 ;
        RECT 2.830000 4.860000 4.030000 5.340000 ;
        RECT 2.830000 10.300000 4.030000 10.780000 ;
        RECT 7.060000 4.860000 8.260000 5.340000 ;
        RECT 7.060000 10.300000 8.260000 10.780000 ;
        RECT 2.830000 15.740000 4.030000 16.220000 ;
        RECT 7.060000 15.740000 8.260000 16.220000 ;
        RECT 2.830000 21.180000 4.030000 21.660000 ;
        RECT 7.060000 21.180000 8.260000 21.660000 ;
        RECT 2.830000 37.500000 4.030000 37.980000 ;
        RECT 7.060000 37.500000 8.260000 37.980000 ;
        RECT 2.830000 26.620000 4.030000 27.100000 ;
        RECT 7.060000 26.620000 8.260000 27.100000 ;
        RECT 2.830000 32.060000 4.030000 32.540000 ;
        RECT 7.060000 32.060000 8.260000 32.540000 ;
        RECT 2.830000 42.940000 4.030000 43.420000 ;
        RECT 7.060000 42.940000 8.260000 43.420000 ;
        RECT 2.830000 48.380000 4.030000 48.860000 ;
        RECT 7.060000 48.380000 8.260000 48.860000 ;
        RECT 52.060000 21.180000 53.260000 21.660000 ;
        RECT 52.060000 15.740000 53.260000 16.220000 ;
        RECT 52.060000 10.300000 53.260000 10.780000 ;
        RECT 52.060000 4.860000 53.260000 5.340000 ;
        RECT 97.060000 21.180000 98.260000 21.660000 ;
        RECT 97.060000 15.740000 98.260000 16.220000 ;
        RECT 97.060000 10.300000 98.260000 10.780000 ;
        RECT 97.060000 4.860000 98.260000 5.340000 ;
        RECT 52.060000 26.620000 53.260000 27.100000 ;
        RECT 52.060000 32.060000 53.260000 32.540000 ;
        RECT 52.060000 37.500000 53.260000 37.980000 ;
        RECT 52.060000 42.940000 53.260000 43.420000 ;
        RECT 52.060000 48.380000 53.260000 48.860000 ;
        RECT 97.060000 26.620000 98.260000 27.100000 ;
        RECT 97.060000 32.060000 98.260000 32.540000 ;
        RECT 97.060000 37.500000 98.260000 37.980000 ;
        RECT 97.060000 42.940000 98.260000 43.420000 ;
        RECT 97.060000 48.380000 98.260000 48.860000 ;
        RECT 2.830000 53.820000 4.030000 54.300000 ;
        RECT 7.060000 53.820000 8.260000 54.300000 ;
        RECT 2.830000 59.260000 4.030000 59.740000 ;
        RECT 7.060000 59.260000 8.260000 59.740000 ;
        RECT 2.830000 64.700000 4.030000 65.180000 ;
        RECT 7.060000 64.700000 8.260000 65.180000 ;
        RECT 2.830000 70.140000 4.030000 70.620000 ;
        RECT 7.060000 70.140000 8.260000 70.620000 ;
        RECT 7.060000 81.020000 8.260000 81.500000 ;
        RECT 2.830000 81.020000 4.030000 81.500000 ;
        RECT 2.830000 75.580000 4.030000 76.060000 ;
        RECT 7.060000 75.580000 8.260000 76.060000 ;
        RECT 2.830000 86.460000 4.030000 86.940000 ;
        RECT 7.060000 86.460000 8.260000 86.940000 ;
        RECT 2.830000 91.900000 4.030000 92.380000 ;
        RECT 7.060000 91.900000 8.260000 92.380000 ;
        RECT 2.830000 97.340000 4.030000 97.820000 ;
        RECT 7.060000 97.340000 8.260000 97.820000 ;
        RECT 52.060000 70.140000 53.260000 70.620000 ;
        RECT 52.060000 53.820000 53.260000 54.300000 ;
        RECT 52.060000 59.260000 53.260000 59.740000 ;
        RECT 52.060000 64.700000 53.260000 65.180000 ;
        RECT 97.060000 53.820000 98.260000 54.300000 ;
        RECT 97.060000 59.260000 98.260000 59.740000 ;
        RECT 97.060000 64.700000 98.260000 65.180000 ;
        RECT 97.060000 70.140000 98.260000 70.620000 ;
        RECT 52.060000 75.580000 53.260000 76.060000 ;
        RECT 52.060000 81.020000 53.260000 81.500000 ;
        RECT 52.060000 86.460000 53.260000 86.940000 ;
        RECT 52.060000 91.900000 53.260000 92.380000 ;
        RECT 52.060000 97.340000 53.260000 97.820000 ;
        RECT 97.060000 75.580000 98.260000 76.060000 ;
        RECT 97.060000 81.020000 98.260000 81.500000 ;
        RECT 97.060000 86.460000 98.260000 86.940000 ;
        RECT 97.060000 91.900000 98.260000 92.380000 ;
        RECT 97.060000 97.340000 98.260000 97.820000 ;
        RECT 142.060000 4.860000 143.260000 5.340000 ;
        RECT 142.060000 10.300000 143.260000 10.780000 ;
        RECT 142.060000 15.740000 143.260000 16.220000 ;
        RECT 142.060000 21.180000 143.260000 21.660000 ;
        RECT 142.060000 26.620000 143.260000 27.100000 ;
        RECT 142.060000 32.060000 143.260000 32.540000 ;
        RECT 142.060000 37.500000 143.260000 37.980000 ;
        RECT 142.060000 42.940000 143.260000 43.420000 ;
        RECT 142.060000 48.380000 143.260000 48.860000 ;
        RECT 196.070000 4.860000 197.270000 5.340000 ;
        RECT 196.070000 10.300000 197.270000 10.780000 ;
        RECT 187.060000 4.860000 188.260000 5.340000 ;
        RECT 187.060000 10.300000 188.260000 10.780000 ;
        RECT 187.060000 15.740000 188.260000 16.220000 ;
        RECT 187.060000 21.180000 188.260000 21.660000 ;
        RECT 196.070000 21.180000 197.270000 21.660000 ;
        RECT 196.070000 15.740000 197.270000 16.220000 ;
        RECT 196.070000 37.500000 197.270000 37.980000 ;
        RECT 187.060000 37.500000 188.260000 37.980000 ;
        RECT 196.070000 26.620000 197.270000 27.100000 ;
        RECT 196.070000 32.060000 197.270000 32.540000 ;
        RECT 187.060000 26.620000 188.260000 27.100000 ;
        RECT 187.060000 32.060000 188.260000 32.540000 ;
        RECT 196.070000 42.940000 197.270000 43.420000 ;
        RECT 196.070000 48.380000 197.270000 48.860000 ;
        RECT 187.060000 42.940000 188.260000 43.420000 ;
        RECT 187.060000 48.380000 188.260000 48.860000 ;
        RECT 142.060000 70.140000 143.260000 70.620000 ;
        RECT 142.060000 64.700000 143.260000 65.180000 ;
        RECT 142.060000 59.260000 143.260000 59.740000 ;
        RECT 142.060000 53.820000 143.260000 54.300000 ;
        RECT 142.060000 75.580000 143.260000 76.060000 ;
        RECT 142.060000 81.020000 143.260000 81.500000 ;
        RECT 142.060000 86.460000 143.260000 86.940000 ;
        RECT 142.060000 91.900000 143.260000 92.380000 ;
        RECT 142.060000 97.340000 143.260000 97.820000 ;
        RECT 187.060000 59.260000 188.260000 59.740000 ;
        RECT 187.060000 53.820000 188.260000 54.300000 ;
        RECT 196.070000 59.260000 197.270000 59.740000 ;
        RECT 196.070000 53.820000 197.270000 54.300000 ;
        RECT 196.070000 64.700000 197.270000 65.180000 ;
        RECT 196.070000 70.140000 197.270000 70.620000 ;
        RECT 187.060000 70.140000 188.260000 70.620000 ;
        RECT 187.060000 64.700000 188.260000 65.180000 ;
        RECT 187.060000 75.580000 188.260000 76.060000 ;
        RECT 187.060000 81.020000 188.260000 81.500000 ;
        RECT 187.060000 86.460000 188.260000 86.940000 ;
        RECT 196.070000 86.460000 197.270000 86.940000 ;
        RECT 196.070000 81.020000 197.270000 81.500000 ;
        RECT 196.070000 75.580000 197.270000 76.060000 ;
        RECT 196.070000 91.900000 197.270000 92.380000 ;
        RECT 196.070000 97.340000 197.270000 97.820000 ;
        RECT 187.060000 91.900000 188.260000 92.380000 ;
        RECT 187.060000 97.340000 188.260000 97.820000 ;
        RECT 2.830000 102.780000 4.030000 103.260000 ;
        RECT 7.060000 102.780000 8.260000 103.260000 ;
        RECT 2.830000 108.220000 4.030000 108.700000 ;
        RECT 7.060000 108.220000 8.260000 108.700000 ;
        RECT 2.830000 113.660000 4.030000 114.140000 ;
        RECT 7.060000 113.660000 8.260000 114.140000 ;
        RECT 2.830000 119.100000 4.030000 119.580000 ;
        RECT 2.830000 124.540000 4.030000 125.020000 ;
        RECT 7.060000 119.100000 8.260000 119.580000 ;
        RECT 7.060000 124.540000 8.260000 125.020000 ;
        RECT 2.830000 129.980000 4.030000 130.460000 ;
        RECT 7.060000 129.980000 8.260000 130.460000 ;
        RECT 2.830000 135.420000 4.030000 135.900000 ;
        RECT 7.060000 135.420000 8.260000 135.900000 ;
        RECT 2.830000 140.860000 4.030000 141.340000 ;
        RECT 7.060000 140.860000 8.260000 141.340000 ;
        RECT 2.830000 146.300000 4.030000 146.780000 ;
        RECT 7.060000 146.300000 8.260000 146.780000 ;
        RECT 52.060000 124.540000 53.260000 125.020000 ;
        RECT 52.060000 119.100000 53.260000 119.580000 ;
        RECT 52.060000 113.660000 53.260000 114.140000 ;
        RECT 52.060000 108.220000 53.260000 108.700000 ;
        RECT 52.060000 102.780000 53.260000 103.260000 ;
        RECT 97.060000 124.540000 98.260000 125.020000 ;
        RECT 97.060000 113.660000 98.260000 114.140000 ;
        RECT 97.060000 108.220000 98.260000 108.700000 ;
        RECT 97.060000 102.780000 98.260000 103.260000 ;
        RECT 97.060000 119.100000 98.260000 119.580000 ;
        RECT 52.060000 129.980000 53.260000 130.460000 ;
        RECT 52.060000 135.420000 53.260000 135.900000 ;
        RECT 52.060000 140.860000 53.260000 141.340000 ;
        RECT 52.060000 146.300000 53.260000 146.780000 ;
        RECT 97.060000 129.980000 98.260000 130.460000 ;
        RECT 97.060000 135.420000 98.260000 135.900000 ;
        RECT 97.060000 140.860000 98.260000 141.340000 ;
        RECT 97.060000 146.300000 98.260000 146.780000 ;
        RECT 2.830000 162.620000 4.030000 163.100000 ;
        RECT 7.060000 162.620000 8.260000 163.100000 ;
        RECT 2.830000 151.740000 4.030000 152.220000 ;
        RECT 7.060000 151.740000 8.260000 152.220000 ;
        RECT 2.830000 157.180000 4.030000 157.660000 ;
        RECT 7.060000 157.180000 8.260000 157.660000 ;
        RECT 2.830000 168.060000 4.030000 168.540000 ;
        RECT 7.060000 168.060000 8.260000 168.540000 ;
        RECT 2.830000 173.500000 4.030000 173.980000 ;
        RECT 7.060000 173.500000 8.260000 173.980000 ;
        RECT 2.830000 178.940000 4.030000 179.420000 ;
        RECT 7.060000 178.940000 8.260000 179.420000 ;
        RECT 7.060000 184.380000 8.260000 184.860000 ;
        RECT 2.830000 184.380000 4.030000 184.860000 ;
        RECT 2.830000 189.820000 4.030000 190.300000 ;
        RECT 7.060000 189.820000 8.260000 190.300000 ;
        RECT 52.060000 168.060000 53.260000 168.540000 ;
        RECT 52.060000 151.740000 53.260000 152.220000 ;
        RECT 52.060000 157.180000 53.260000 157.660000 ;
        RECT 52.060000 162.620000 53.260000 163.100000 ;
        RECT 52.060000 173.500000 53.260000 173.980000 ;
        RECT 97.060000 173.500000 98.260000 173.980000 ;
        RECT 97.060000 168.060000 98.260000 168.540000 ;
        RECT 97.060000 151.740000 98.260000 152.220000 ;
        RECT 97.060000 157.180000 98.260000 157.660000 ;
        RECT 97.060000 162.620000 98.260000 163.100000 ;
        RECT 52.060000 178.940000 53.260000 179.420000 ;
        RECT 52.060000 184.380000 53.260000 184.860000 ;
        RECT 52.060000 189.820000 53.260000 190.300000 ;
        RECT 97.060000 178.940000 98.260000 179.420000 ;
        RECT 97.060000 184.380000 98.260000 184.860000 ;
        RECT 97.060000 189.820000 98.260000 190.300000 ;
        RECT 142.060000 124.540000 143.260000 125.020000 ;
        RECT 142.060000 102.780000 143.260000 103.260000 ;
        RECT 142.060000 108.220000 143.260000 108.700000 ;
        RECT 142.060000 113.660000 143.260000 114.140000 ;
        RECT 142.060000 119.100000 143.260000 119.580000 ;
        RECT 142.060000 129.980000 143.260000 130.460000 ;
        RECT 142.060000 135.420000 143.260000 135.900000 ;
        RECT 142.060000 140.860000 143.260000 141.340000 ;
        RECT 142.060000 146.300000 143.260000 146.780000 ;
        RECT 196.070000 102.780000 197.270000 103.260000 ;
        RECT 196.070000 108.220000 197.270000 108.700000 ;
        RECT 187.060000 102.780000 188.260000 103.260000 ;
        RECT 187.060000 108.220000 188.260000 108.700000 ;
        RECT 187.060000 124.540000 188.260000 125.020000 ;
        RECT 187.060000 113.660000 188.260000 114.140000 ;
        RECT 187.060000 119.100000 188.260000 119.580000 ;
        RECT 196.070000 124.540000 197.270000 125.020000 ;
        RECT 196.070000 119.100000 197.270000 119.580000 ;
        RECT 196.070000 113.660000 197.270000 114.140000 ;
        RECT 196.070000 129.980000 197.270000 130.460000 ;
        RECT 196.070000 135.420000 197.270000 135.900000 ;
        RECT 187.060000 129.980000 188.260000 130.460000 ;
        RECT 187.060000 135.420000 188.260000 135.900000 ;
        RECT 187.060000 140.860000 188.260000 141.340000 ;
        RECT 187.060000 146.300000 188.260000 146.780000 ;
        RECT 196.070000 146.300000 197.270000 146.780000 ;
        RECT 196.070000 140.860000 197.270000 141.340000 ;
        RECT 142.060000 168.060000 143.260000 168.540000 ;
        RECT 142.060000 162.620000 143.260000 163.100000 ;
        RECT 142.060000 157.180000 143.260000 157.660000 ;
        RECT 142.060000 151.740000 143.260000 152.220000 ;
        RECT 142.060000 173.500000 143.260000 173.980000 ;
        RECT 142.060000 178.940000 143.260000 179.420000 ;
        RECT 142.060000 184.380000 143.260000 184.860000 ;
        RECT 142.060000 189.820000 143.260000 190.300000 ;
        RECT 196.070000 162.620000 197.270000 163.100000 ;
        RECT 187.060000 162.620000 188.260000 163.100000 ;
        RECT 196.070000 151.740000 197.270000 152.220000 ;
        RECT 196.070000 157.180000 197.270000 157.660000 ;
        RECT 187.060000 157.180000 188.260000 157.660000 ;
        RECT 187.060000 151.740000 188.260000 152.220000 ;
        RECT 196.070000 168.060000 197.270000 168.540000 ;
        RECT 196.070000 173.500000 197.270000 173.980000 ;
        RECT 187.060000 168.060000 188.260000 168.540000 ;
        RECT 187.060000 173.500000 188.260000 173.980000 ;
        RECT 187.060000 178.940000 188.260000 179.420000 ;
        RECT 187.060000 184.380000 188.260000 184.860000 ;
        RECT 196.070000 184.380000 197.270000 184.860000 ;
        RECT 196.070000 178.940000 197.270000 179.420000 ;
        RECT 196.070000 189.820000 197.270000 190.300000 ;
        RECT 187.060000 189.820000 188.260000 190.300000 ;
      LAYER met4 ;
        RECT 2.830000 0.000000 4.030000 200.260000 ;
        RECT 7.060000 2.850000 8.260000 196.220000 ;
        RECT 52.060000 2.850000 53.260000 196.220000 ;
        RECT 97.060000 2.850000 98.260000 196.220000 ;
        RECT 196.070000 0.000000 197.270000 200.260000 ;
        RECT 142.060000 2.850000 143.260000 196.220000 ;
        RECT 187.060000 2.850000 188.260000 196.220000 ;
    END
# end of P/G power stripe data as pin

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 198.900000 196.820000 200.100000 198.020000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 196.820000 1.200000 198.020000 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.900000 1.050000 200.100000 2.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 1.200000 2.250000 ;
    END
    PORT
      LAYER met4 ;
        RECT 197.870000 199.060000 199.070000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 197.870000 0.000000 199.070000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 199.060000 2.230000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 0.000000 2.230000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 200.100000 2.250000 ;
        RECT 0.000000 196.820000 200.100000 198.020000 ;
        RECT 4.895000 100.060000 6.260000 100.540000 ;
        RECT 1.030000 100.060000 2.230000 100.540000 ;
        RECT 95.060000 100.060000 96.260000 100.540000 ;
        RECT 50.060000 100.060000 51.260000 100.540000 ;
        RECT 197.870000 100.060000 199.070000 100.540000 ;
        RECT 185.060000 100.060000 186.260000 100.540000 ;
        RECT 140.060000 100.060000 141.260000 100.540000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 1.030000 7.580000 2.230000 8.060000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 1.030000 18.460000 2.230000 18.940000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 1.030000 13.020000 2.230000 13.500000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
        RECT 1.030000 23.900000 2.230000 24.380000 ;
        RECT 4.895000 29.340000 6.260000 29.820000 ;
        RECT 1.030000 29.340000 2.230000 29.820000 ;
        RECT 4.895000 34.780000 6.260000 35.260000 ;
        RECT 1.030000 34.780000 2.230000 35.260000 ;
        RECT 4.895000 40.220000 6.260000 40.700000 ;
        RECT 1.030000 40.220000 2.230000 40.700000 ;
        RECT 4.895000 45.660000 6.260000 46.140000 ;
        RECT 1.030000 45.660000 2.230000 46.140000 ;
        RECT 50.060000 23.900000 51.260000 24.380000 ;
        RECT 50.060000 18.460000 51.260000 18.940000 ;
        RECT 50.060000 13.020000 51.260000 13.500000 ;
        RECT 50.060000 7.580000 51.260000 8.060000 ;
        RECT 95.060000 23.900000 96.260000 24.380000 ;
        RECT 95.060000 18.460000 96.260000 18.940000 ;
        RECT 95.060000 13.020000 96.260000 13.500000 ;
        RECT 95.060000 7.580000 96.260000 8.060000 ;
        RECT 50.060000 45.660000 51.260000 46.140000 ;
        RECT 50.060000 40.220000 51.260000 40.700000 ;
        RECT 50.060000 34.780000 51.260000 35.260000 ;
        RECT 50.060000 29.340000 51.260000 29.820000 ;
        RECT 95.060000 45.660000 96.260000 46.140000 ;
        RECT 95.060000 40.220000 96.260000 40.700000 ;
        RECT 95.060000 34.780000 96.260000 35.260000 ;
        RECT 95.060000 29.340000 96.260000 29.820000 ;
        RECT 4.895000 51.100000 6.260000 51.580000 ;
        RECT 1.030000 51.100000 2.230000 51.580000 ;
        RECT 4.895000 61.980000 6.260000 62.460000 ;
        RECT 1.030000 61.980000 2.230000 62.460000 ;
        RECT 4.895000 56.540000 6.260000 57.020000 ;
        RECT 1.030000 56.540000 2.230000 57.020000 ;
        RECT 4.895000 67.420000 6.260000 67.900000 ;
        RECT 1.030000 67.420000 2.230000 67.900000 ;
        RECT 4.895000 72.860000 6.260000 73.340000 ;
        RECT 1.030000 72.860000 2.230000 73.340000 ;
        RECT 4.895000 78.300000 6.260000 78.780000 ;
        RECT 1.030000 78.300000 2.230000 78.780000 ;
        RECT 4.895000 83.740000 6.260000 84.220000 ;
        RECT 1.030000 83.740000 2.230000 84.220000 ;
        RECT 4.895000 89.180000 6.260000 89.660000 ;
        RECT 1.030000 89.180000 2.230000 89.660000 ;
        RECT 4.895000 94.620000 6.260000 95.100000 ;
        RECT 1.030000 94.620000 2.230000 95.100000 ;
        RECT 50.060000 72.860000 51.260000 73.340000 ;
        RECT 50.060000 67.420000 51.260000 67.900000 ;
        RECT 50.060000 61.980000 51.260000 62.460000 ;
        RECT 50.060000 56.540000 51.260000 57.020000 ;
        RECT 50.060000 51.100000 51.260000 51.580000 ;
        RECT 95.060000 72.860000 96.260000 73.340000 ;
        RECT 95.060000 67.420000 96.260000 67.900000 ;
        RECT 95.060000 61.980000 96.260000 62.460000 ;
        RECT 95.060000 56.540000 96.260000 57.020000 ;
        RECT 95.060000 51.100000 96.260000 51.580000 ;
        RECT 50.060000 94.620000 51.260000 95.100000 ;
        RECT 50.060000 89.180000 51.260000 89.660000 ;
        RECT 50.060000 83.740000 51.260000 84.220000 ;
        RECT 50.060000 78.300000 51.260000 78.780000 ;
        RECT 95.060000 94.620000 96.260000 95.100000 ;
        RECT 95.060000 89.180000 96.260000 89.660000 ;
        RECT 95.060000 83.740000 96.260000 84.220000 ;
        RECT 95.060000 78.300000 96.260000 78.780000 ;
        RECT 140.060000 23.900000 141.260000 24.380000 ;
        RECT 140.060000 18.460000 141.260000 18.940000 ;
        RECT 140.060000 13.020000 141.260000 13.500000 ;
        RECT 140.060000 7.580000 141.260000 8.060000 ;
        RECT 140.060000 45.660000 141.260000 46.140000 ;
        RECT 140.060000 40.220000 141.260000 40.700000 ;
        RECT 140.060000 34.780000 141.260000 35.260000 ;
        RECT 140.060000 29.340000 141.260000 29.820000 ;
        RECT 197.870000 7.580000 199.070000 8.060000 ;
        RECT 185.060000 7.580000 186.260000 8.060000 ;
        RECT 185.060000 13.020000 186.260000 13.500000 ;
        RECT 185.060000 18.460000 186.260000 18.940000 ;
        RECT 185.060000 23.900000 186.260000 24.380000 ;
        RECT 197.870000 23.900000 199.070000 24.380000 ;
        RECT 197.870000 13.020000 199.070000 13.500000 ;
        RECT 197.870000 18.460000 199.070000 18.940000 ;
        RECT 197.870000 34.780000 199.070000 35.260000 ;
        RECT 197.870000 29.340000 199.070000 29.820000 ;
        RECT 185.060000 34.780000 186.260000 35.260000 ;
        RECT 185.060000 29.340000 186.260000 29.820000 ;
        RECT 197.870000 45.660000 199.070000 46.140000 ;
        RECT 197.870000 40.220000 199.070000 40.700000 ;
        RECT 185.060000 45.660000 186.260000 46.140000 ;
        RECT 185.060000 40.220000 186.260000 40.700000 ;
        RECT 140.060000 72.860000 141.260000 73.340000 ;
        RECT 140.060000 67.420000 141.260000 67.900000 ;
        RECT 140.060000 61.980000 141.260000 62.460000 ;
        RECT 140.060000 56.540000 141.260000 57.020000 ;
        RECT 140.060000 51.100000 141.260000 51.580000 ;
        RECT 140.060000 94.620000 141.260000 95.100000 ;
        RECT 140.060000 89.180000 141.260000 89.660000 ;
        RECT 140.060000 83.740000 141.260000 84.220000 ;
        RECT 140.060000 78.300000 141.260000 78.780000 ;
        RECT 185.060000 51.100000 186.260000 51.580000 ;
        RECT 185.060000 56.540000 186.260000 57.020000 ;
        RECT 185.060000 61.980000 186.260000 62.460000 ;
        RECT 197.870000 61.980000 199.070000 62.460000 ;
        RECT 197.870000 51.100000 199.070000 51.580000 ;
        RECT 197.870000 56.540000 199.070000 57.020000 ;
        RECT 197.870000 72.860000 199.070000 73.340000 ;
        RECT 197.870000 67.420000 199.070000 67.900000 ;
        RECT 185.060000 72.860000 186.260000 73.340000 ;
        RECT 185.060000 67.420000 186.260000 67.900000 ;
        RECT 185.060000 78.300000 186.260000 78.780000 ;
        RECT 185.060000 83.740000 186.260000 84.220000 ;
        RECT 197.870000 83.740000 199.070000 84.220000 ;
        RECT 197.870000 78.300000 199.070000 78.780000 ;
        RECT 197.870000 94.620000 199.070000 95.100000 ;
        RECT 197.870000 89.180000 199.070000 89.660000 ;
        RECT 185.060000 94.620000 186.260000 95.100000 ;
        RECT 185.060000 89.180000 186.260000 89.660000 ;
        RECT 4.895000 105.500000 6.260000 105.980000 ;
        RECT 1.030000 105.500000 2.230000 105.980000 ;
        RECT 4.895000 110.940000 6.260000 111.420000 ;
        RECT 1.030000 110.940000 2.230000 111.420000 ;
        RECT 4.895000 116.380000 6.260000 116.860000 ;
        RECT 1.030000 116.380000 2.230000 116.860000 ;
        RECT 4.895000 121.820000 6.260000 122.300000 ;
        RECT 1.030000 121.820000 2.230000 122.300000 ;
        RECT 4.895000 127.260000 6.260000 127.740000 ;
        RECT 1.030000 127.260000 2.230000 127.740000 ;
        RECT 4.895000 132.700000 6.260000 133.180000 ;
        RECT 1.030000 132.700000 2.230000 133.180000 ;
        RECT 4.895000 143.580000 6.260000 144.060000 ;
        RECT 1.030000 143.580000 2.230000 144.060000 ;
        RECT 4.895000 138.140000 6.260000 138.620000 ;
        RECT 1.030000 138.140000 2.230000 138.620000 ;
        RECT 4.895000 149.020000 6.260000 149.500000 ;
        RECT 1.030000 149.020000 2.230000 149.500000 ;
        RECT 50.060000 121.820000 51.260000 122.300000 ;
        RECT 50.060000 116.380000 51.260000 116.860000 ;
        RECT 50.060000 110.940000 51.260000 111.420000 ;
        RECT 50.060000 105.500000 51.260000 105.980000 ;
        RECT 95.060000 121.820000 96.260000 122.300000 ;
        RECT 95.060000 116.380000 96.260000 116.860000 ;
        RECT 95.060000 110.940000 96.260000 111.420000 ;
        RECT 95.060000 105.500000 96.260000 105.980000 ;
        RECT 50.060000 149.020000 51.260000 149.500000 ;
        RECT 50.060000 143.580000 51.260000 144.060000 ;
        RECT 50.060000 138.140000 51.260000 138.620000 ;
        RECT 50.060000 132.700000 51.260000 133.180000 ;
        RECT 50.060000 127.260000 51.260000 127.740000 ;
        RECT 95.060000 149.020000 96.260000 149.500000 ;
        RECT 95.060000 143.580000 96.260000 144.060000 ;
        RECT 95.060000 138.140000 96.260000 138.620000 ;
        RECT 95.060000 132.700000 96.260000 133.180000 ;
        RECT 95.060000 127.260000 96.260000 127.740000 ;
        RECT 4.895000 154.460000 6.260000 154.940000 ;
        RECT 1.030000 154.460000 2.230000 154.940000 ;
        RECT 4.895000 159.900000 6.260000 160.380000 ;
        RECT 1.030000 159.900000 2.230000 160.380000 ;
        RECT 4.895000 165.340000 6.260000 165.820000 ;
        RECT 1.030000 165.340000 2.230000 165.820000 ;
        RECT 4.895000 170.780000 6.260000 171.260000 ;
        RECT 1.030000 170.780000 2.230000 171.260000 ;
        RECT 4.895000 176.220000 6.260000 176.700000 ;
        RECT 1.030000 176.220000 2.230000 176.700000 ;
        RECT 4.895000 187.100000 6.260000 187.580000 ;
        RECT 1.030000 187.100000 2.230000 187.580000 ;
        RECT 4.895000 181.660000 6.260000 182.140000 ;
        RECT 1.030000 181.660000 2.230000 182.140000 ;
        RECT 4.895000 192.540000 6.260000 193.020000 ;
        RECT 1.030000 192.540000 2.230000 193.020000 ;
        RECT 50.060000 170.780000 51.260000 171.260000 ;
        RECT 50.060000 165.340000 51.260000 165.820000 ;
        RECT 50.060000 159.900000 51.260000 160.380000 ;
        RECT 50.060000 154.460000 51.260000 154.940000 ;
        RECT 95.060000 170.780000 96.260000 171.260000 ;
        RECT 95.060000 165.340000 96.260000 165.820000 ;
        RECT 95.060000 159.900000 96.260000 160.380000 ;
        RECT 95.060000 154.460000 96.260000 154.940000 ;
        RECT 50.060000 192.540000 51.260000 193.020000 ;
        RECT 50.060000 187.100000 51.260000 187.580000 ;
        RECT 50.060000 181.660000 51.260000 182.140000 ;
        RECT 50.060000 176.220000 51.260000 176.700000 ;
        RECT 95.060000 192.540000 96.260000 193.020000 ;
        RECT 95.060000 187.100000 96.260000 187.580000 ;
        RECT 95.060000 176.220000 96.260000 176.700000 ;
        RECT 95.060000 181.660000 96.260000 182.140000 ;
        RECT 140.060000 121.820000 141.260000 122.300000 ;
        RECT 140.060000 116.380000 141.260000 116.860000 ;
        RECT 140.060000 110.940000 141.260000 111.420000 ;
        RECT 140.060000 105.500000 141.260000 105.980000 ;
        RECT 140.060000 149.020000 141.260000 149.500000 ;
        RECT 140.060000 143.580000 141.260000 144.060000 ;
        RECT 140.060000 138.140000 141.260000 138.620000 ;
        RECT 140.060000 132.700000 141.260000 133.180000 ;
        RECT 140.060000 127.260000 141.260000 127.740000 ;
        RECT 197.870000 110.940000 199.070000 111.420000 ;
        RECT 197.870000 105.500000 199.070000 105.980000 ;
        RECT 185.060000 110.940000 186.260000 111.420000 ;
        RECT 185.060000 105.500000 186.260000 105.980000 ;
        RECT 185.060000 116.380000 186.260000 116.860000 ;
        RECT 185.060000 121.820000 186.260000 122.300000 ;
        RECT 197.870000 121.820000 199.070000 122.300000 ;
        RECT 197.870000 116.380000 199.070000 116.860000 ;
        RECT 197.870000 132.700000 199.070000 133.180000 ;
        RECT 197.870000 127.260000 199.070000 127.740000 ;
        RECT 185.060000 132.700000 186.260000 133.180000 ;
        RECT 185.060000 127.260000 186.260000 127.740000 ;
        RECT 185.060000 138.140000 186.260000 138.620000 ;
        RECT 185.060000 143.580000 186.260000 144.060000 ;
        RECT 185.060000 149.020000 186.260000 149.500000 ;
        RECT 197.870000 149.020000 199.070000 149.500000 ;
        RECT 197.870000 138.140000 199.070000 138.620000 ;
        RECT 197.870000 143.580000 199.070000 144.060000 ;
        RECT 140.060000 170.780000 141.260000 171.260000 ;
        RECT 140.060000 165.340000 141.260000 165.820000 ;
        RECT 140.060000 154.460000 141.260000 154.940000 ;
        RECT 140.060000 159.900000 141.260000 160.380000 ;
        RECT 140.060000 192.540000 141.260000 193.020000 ;
        RECT 140.060000 187.100000 141.260000 187.580000 ;
        RECT 140.060000 181.660000 141.260000 182.140000 ;
        RECT 140.060000 176.220000 141.260000 176.700000 ;
        RECT 197.870000 159.900000 199.070000 160.380000 ;
        RECT 197.870000 154.460000 199.070000 154.940000 ;
        RECT 185.060000 159.900000 186.260000 160.380000 ;
        RECT 185.060000 154.460000 186.260000 154.940000 ;
        RECT 197.870000 170.780000 199.070000 171.260000 ;
        RECT 197.870000 165.340000 199.070000 165.820000 ;
        RECT 185.060000 170.780000 186.260000 171.260000 ;
        RECT 185.060000 165.340000 186.260000 165.820000 ;
        RECT 185.060000 176.220000 186.260000 176.700000 ;
        RECT 185.060000 181.660000 186.260000 182.140000 ;
        RECT 185.060000 187.100000 186.260000 187.580000 ;
        RECT 197.870000 187.100000 199.070000 187.580000 ;
        RECT 197.870000 176.220000 199.070000 176.700000 ;
        RECT 197.870000 181.660000 199.070000 182.140000 ;
        RECT 197.870000 192.540000 199.070000 193.020000 ;
        RECT 185.060000 192.540000 186.260000 193.020000 ;
      LAYER met4 ;
        RECT 1.030000 0.000000 2.230000 200.260000 ;
        RECT 5.060000 1.050000 6.260000 198.020000 ;
        RECT 50.060000 1.050000 51.260000 198.020000 ;
        RECT 95.060000 1.050000 96.260000 198.020000 ;
        RECT 197.870000 0.000000 199.070000 200.260000 ;
        RECT 140.060000 1.050000 141.260000 198.020000 ;
        RECT 185.060000 1.050000 186.260000 198.020000 ;
        RECT 4.895000 100.060000 6.260000 100.540000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
        RECT 4.895000 29.340000 6.260000 29.820000 ;
        RECT 4.895000 34.780000 6.260000 35.260000 ;
        RECT 4.895000 40.220000 6.260000 40.700000 ;
        RECT 4.895000 45.660000 6.260000 46.140000 ;
        RECT 4.895000 51.100000 6.260000 51.580000 ;
        RECT 4.895000 61.980000 6.260000 62.460000 ;
        RECT 4.895000 56.540000 6.260000 57.020000 ;
        RECT 4.895000 67.420000 6.260000 67.900000 ;
        RECT 4.895000 72.860000 6.260000 73.340000 ;
        RECT 4.895000 78.300000 6.260000 78.780000 ;
        RECT 4.895000 83.740000 6.260000 84.220000 ;
        RECT 4.895000 89.180000 6.260000 89.660000 ;
        RECT 4.895000 94.620000 6.260000 95.100000 ;
        RECT 4.895000 105.500000 6.260000 105.980000 ;
        RECT 4.895000 110.940000 6.260000 111.420000 ;
        RECT 4.895000 116.380000 6.260000 116.860000 ;
        RECT 4.895000 121.820000 6.260000 122.300000 ;
        RECT 4.895000 127.260000 6.260000 127.740000 ;
        RECT 4.895000 132.700000 6.260000 133.180000 ;
        RECT 4.895000 143.580000 6.260000 144.060000 ;
        RECT 4.895000 138.140000 6.260000 138.620000 ;
        RECT 4.895000 149.020000 6.260000 149.500000 ;
        RECT 4.895000 154.460000 6.260000 154.940000 ;
        RECT 4.895000 159.900000 6.260000 160.380000 ;
        RECT 4.895000 165.340000 6.260000 165.820000 ;
        RECT 4.895000 170.780000 6.260000 171.260000 ;
        RECT 4.895000 176.220000 6.260000 176.700000 ;
        RECT 4.895000 187.100000 6.260000 187.580000 ;
        RECT 4.895000 181.660000 6.260000 182.140000 ;
        RECT 4.895000 192.540000 6.260000 193.020000 ;
    END
# end of P/G power stripe data as pin

  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 200.100000 200.260000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 200.100000 200.260000 ;
    LAYER met2 ;
      RECT 194.680000 199.420000 200.100000 200.260000 ;
      RECT 193.300000 199.420000 194.020000 200.260000 ;
      RECT 191.920000 199.420000 192.640000 200.260000 ;
      RECT 190.540000 199.420000 191.260000 200.260000 ;
      RECT 188.700000 199.420000 189.880000 200.260000 ;
      RECT 187.320000 199.420000 188.040000 200.260000 ;
      RECT 185.940000 199.420000 186.660000 200.260000 ;
      RECT 184.100000 199.420000 185.280000 200.260000 ;
      RECT 182.720000 199.420000 183.440000 200.260000 ;
      RECT 181.340000 199.420000 182.060000 200.260000 ;
      RECT 179.960000 199.420000 180.680000 200.260000 ;
      RECT 178.120000 199.420000 179.300000 200.260000 ;
      RECT 176.740000 199.420000 177.460000 200.260000 ;
      RECT 175.360000 199.420000 176.080000 200.260000 ;
      RECT 173.520000 199.420000 174.700000 200.260000 ;
      RECT 172.140000 199.420000 172.860000 200.260000 ;
      RECT 170.760000 199.420000 171.480000 200.260000 ;
      RECT 168.920000 199.420000 170.100000 200.260000 ;
      RECT 167.540000 199.420000 168.260000 200.260000 ;
      RECT 166.160000 199.420000 166.880000 200.260000 ;
      RECT 164.780000 199.420000 165.500000 200.260000 ;
      RECT 162.940000 199.420000 164.120000 200.260000 ;
      RECT 161.560000 199.420000 162.280000 200.260000 ;
      RECT 160.180000 199.420000 160.900000 200.260000 ;
      RECT 158.340000 199.420000 159.520000 200.260000 ;
      RECT 156.960000 199.420000 157.680000 200.260000 ;
      RECT 155.580000 199.420000 156.300000 200.260000 ;
      RECT 154.200000 199.420000 154.920000 200.260000 ;
      RECT 152.360000 199.420000 153.540000 200.260000 ;
      RECT 150.980000 199.420000 151.700000 200.260000 ;
      RECT 149.600000 199.420000 150.320000 200.260000 ;
      RECT 147.760000 199.420000 148.940000 200.260000 ;
      RECT 146.380000 199.420000 147.100000 200.260000 ;
      RECT 145.000000 199.420000 145.720000 200.260000 ;
      RECT 143.160000 199.420000 144.340000 200.260000 ;
      RECT 141.780000 199.420000 142.500000 200.260000 ;
      RECT 140.400000 199.420000 141.120000 200.260000 ;
      RECT 139.020000 199.420000 139.740000 200.260000 ;
      RECT 137.180000 199.420000 138.360000 200.260000 ;
      RECT 135.800000 199.420000 136.520000 200.260000 ;
      RECT 134.420000 199.420000 135.140000 200.260000 ;
      RECT 132.580000 199.420000 133.760000 200.260000 ;
      RECT 131.200000 199.420000 131.920000 200.260000 ;
      RECT 129.820000 199.420000 130.540000 200.260000 ;
      RECT 127.980000 199.420000 129.160000 200.260000 ;
      RECT 126.600000 199.420000 127.320000 200.260000 ;
      RECT 125.220000 199.420000 125.940000 200.260000 ;
      RECT 123.840000 199.420000 124.560000 200.260000 ;
      RECT 122.000000 199.420000 123.180000 200.260000 ;
      RECT 120.620000 199.420000 121.340000 200.260000 ;
      RECT 119.240000 199.420000 119.960000 200.260000 ;
      RECT 117.400000 199.420000 118.580000 200.260000 ;
      RECT 116.020000 199.420000 116.740000 200.260000 ;
      RECT 114.640000 199.420000 115.360000 200.260000 ;
      RECT 113.260000 199.420000 113.980000 200.260000 ;
      RECT 111.420000 199.420000 112.600000 200.260000 ;
      RECT 110.040000 199.420000 110.760000 200.260000 ;
      RECT 108.660000 199.420000 109.380000 200.260000 ;
      RECT 106.820000 199.420000 108.000000 200.260000 ;
      RECT 105.440000 199.420000 106.160000 200.260000 ;
      RECT 104.060000 199.420000 104.780000 200.260000 ;
      RECT 102.220000 199.420000 103.400000 200.260000 ;
      RECT 100.840000 199.420000 101.560000 200.260000 ;
      RECT 99.460000 199.420000 100.180000 200.260000 ;
      RECT 98.080000 199.420000 98.800000 200.260000 ;
      RECT 96.240000 199.420000 97.420000 200.260000 ;
      RECT 94.860000 199.420000 95.580000 200.260000 ;
      RECT 93.480000 199.420000 94.200000 200.260000 ;
      RECT 91.640000 199.420000 92.820000 200.260000 ;
      RECT 90.260000 199.420000 90.980000 200.260000 ;
      RECT 88.880000 199.420000 89.600000 200.260000 ;
      RECT 87.040000 199.420000 88.220000 200.260000 ;
      RECT 85.660000 199.420000 86.380000 200.260000 ;
      RECT 84.280000 199.420000 85.000000 200.260000 ;
      RECT 82.900000 199.420000 83.620000 200.260000 ;
      RECT 81.060000 199.420000 82.240000 200.260000 ;
      RECT 79.680000 199.420000 80.400000 200.260000 ;
      RECT 78.300000 199.420000 79.020000 200.260000 ;
      RECT 76.460000 199.420000 77.640000 200.260000 ;
      RECT 75.080000 199.420000 75.800000 200.260000 ;
      RECT 73.700000 199.420000 74.420000 200.260000 ;
      RECT 72.320000 199.420000 73.040000 200.260000 ;
      RECT 70.480000 199.420000 71.660000 200.260000 ;
      RECT 69.100000 199.420000 69.820000 200.260000 ;
      RECT 67.720000 199.420000 68.440000 200.260000 ;
      RECT 65.880000 199.420000 67.060000 200.260000 ;
      RECT 64.500000 199.420000 65.220000 200.260000 ;
      RECT 63.120000 199.420000 63.840000 200.260000 ;
      RECT 61.280000 199.420000 62.460000 200.260000 ;
      RECT 59.900000 199.420000 60.620000 200.260000 ;
      RECT 58.520000 199.420000 59.240000 200.260000 ;
      RECT 57.140000 199.420000 57.860000 200.260000 ;
      RECT 55.300000 199.420000 56.480000 200.260000 ;
      RECT 53.920000 199.420000 54.640000 200.260000 ;
      RECT 52.540000 199.420000 53.260000 200.260000 ;
      RECT 50.700000 199.420000 51.880000 200.260000 ;
      RECT 49.320000 199.420000 50.040000 200.260000 ;
      RECT 47.940000 199.420000 48.660000 200.260000 ;
      RECT 46.100000 199.420000 47.280000 200.260000 ;
      RECT 44.720000 199.420000 45.440000 200.260000 ;
      RECT 43.340000 199.420000 44.060000 200.260000 ;
      RECT 41.960000 199.420000 42.680000 200.260000 ;
      RECT 40.120000 199.420000 41.300000 200.260000 ;
      RECT 38.740000 199.420000 39.460000 200.260000 ;
      RECT 37.360000 199.420000 38.080000 200.260000 ;
      RECT 35.520000 199.420000 36.700000 200.260000 ;
      RECT 34.140000 199.420000 34.860000 200.260000 ;
      RECT 32.760000 199.420000 33.480000 200.260000 ;
      RECT 31.380000 199.420000 32.100000 200.260000 ;
      RECT 29.540000 199.420000 30.720000 200.260000 ;
      RECT 28.160000 199.420000 28.880000 200.260000 ;
      RECT 26.780000 199.420000 27.500000 200.260000 ;
      RECT 24.940000 199.420000 26.120000 200.260000 ;
      RECT 23.560000 199.420000 24.280000 200.260000 ;
      RECT 22.180000 199.420000 22.900000 200.260000 ;
      RECT 20.340000 199.420000 21.520000 200.260000 ;
      RECT 18.960000 199.420000 19.680000 200.260000 ;
      RECT 17.580000 199.420000 18.300000 200.260000 ;
      RECT 16.200000 199.420000 16.920000 200.260000 ;
      RECT 14.360000 199.420000 15.540000 200.260000 ;
      RECT 12.980000 199.420000 13.700000 200.260000 ;
      RECT 11.600000 199.420000 12.320000 200.260000 ;
      RECT 9.760000 199.420000 10.940000 200.260000 ;
      RECT 8.380000 199.420000 9.100000 200.260000 ;
      RECT 7.000000 199.420000 7.720000 200.260000 ;
      RECT 5.620000 199.420000 6.340000 200.260000 ;
      RECT 0.000000 199.420000 4.960000 200.260000 ;
      RECT 0.000000 0.840000 200.100000 199.420000 ;
      RECT 194.680000 0.000000 200.100000 0.840000 ;
      RECT 193.300000 0.000000 194.020000 0.840000 ;
      RECT 191.920000 0.000000 192.640000 0.840000 ;
      RECT 190.540000 0.000000 191.260000 0.840000 ;
      RECT 188.700000 0.000000 189.880000 0.840000 ;
      RECT 187.320000 0.000000 188.040000 0.840000 ;
      RECT 185.940000 0.000000 186.660000 0.840000 ;
      RECT 184.100000 0.000000 185.280000 0.840000 ;
      RECT 182.720000 0.000000 183.440000 0.840000 ;
      RECT 181.340000 0.000000 182.060000 0.840000 ;
      RECT 179.960000 0.000000 180.680000 0.840000 ;
      RECT 178.120000 0.000000 179.300000 0.840000 ;
      RECT 176.740000 0.000000 177.460000 0.840000 ;
      RECT 175.360000 0.000000 176.080000 0.840000 ;
      RECT 173.520000 0.000000 174.700000 0.840000 ;
      RECT 172.140000 0.000000 172.860000 0.840000 ;
      RECT 170.760000 0.000000 171.480000 0.840000 ;
      RECT 168.920000 0.000000 170.100000 0.840000 ;
      RECT 167.540000 0.000000 168.260000 0.840000 ;
      RECT 166.160000 0.000000 166.880000 0.840000 ;
      RECT 164.780000 0.000000 165.500000 0.840000 ;
      RECT 162.940000 0.000000 164.120000 0.840000 ;
      RECT 161.560000 0.000000 162.280000 0.840000 ;
      RECT 160.180000 0.000000 160.900000 0.840000 ;
      RECT 158.340000 0.000000 159.520000 0.840000 ;
      RECT 156.960000 0.000000 157.680000 0.840000 ;
      RECT 155.580000 0.000000 156.300000 0.840000 ;
      RECT 154.200000 0.000000 154.920000 0.840000 ;
      RECT 152.360000 0.000000 153.540000 0.840000 ;
      RECT 150.980000 0.000000 151.700000 0.840000 ;
      RECT 149.600000 0.000000 150.320000 0.840000 ;
      RECT 147.760000 0.000000 148.940000 0.840000 ;
      RECT 146.380000 0.000000 147.100000 0.840000 ;
      RECT 145.000000 0.000000 145.720000 0.840000 ;
      RECT 143.160000 0.000000 144.340000 0.840000 ;
      RECT 141.780000 0.000000 142.500000 0.840000 ;
      RECT 140.400000 0.000000 141.120000 0.840000 ;
      RECT 139.020000 0.000000 139.740000 0.840000 ;
      RECT 137.180000 0.000000 138.360000 0.840000 ;
      RECT 135.800000 0.000000 136.520000 0.840000 ;
      RECT 134.420000 0.000000 135.140000 0.840000 ;
      RECT 132.580000 0.000000 133.760000 0.840000 ;
      RECT 131.200000 0.000000 131.920000 0.840000 ;
      RECT 129.820000 0.000000 130.540000 0.840000 ;
      RECT 127.980000 0.000000 129.160000 0.840000 ;
      RECT 126.600000 0.000000 127.320000 0.840000 ;
      RECT 125.220000 0.000000 125.940000 0.840000 ;
      RECT 123.840000 0.000000 124.560000 0.840000 ;
      RECT 122.000000 0.000000 123.180000 0.840000 ;
      RECT 120.620000 0.000000 121.340000 0.840000 ;
      RECT 119.240000 0.000000 119.960000 0.840000 ;
      RECT 117.400000 0.000000 118.580000 0.840000 ;
      RECT 116.020000 0.000000 116.740000 0.840000 ;
      RECT 114.640000 0.000000 115.360000 0.840000 ;
      RECT 113.260000 0.000000 113.980000 0.840000 ;
      RECT 111.420000 0.000000 112.600000 0.840000 ;
      RECT 110.040000 0.000000 110.760000 0.840000 ;
      RECT 108.660000 0.000000 109.380000 0.840000 ;
      RECT 106.820000 0.000000 108.000000 0.840000 ;
      RECT 105.440000 0.000000 106.160000 0.840000 ;
      RECT 104.060000 0.000000 104.780000 0.840000 ;
      RECT 102.220000 0.000000 103.400000 0.840000 ;
      RECT 100.840000 0.000000 101.560000 0.840000 ;
      RECT 99.460000 0.000000 100.180000 0.840000 ;
      RECT 98.080000 0.000000 98.800000 0.840000 ;
      RECT 96.240000 0.000000 97.420000 0.840000 ;
      RECT 94.860000 0.000000 95.580000 0.840000 ;
      RECT 93.480000 0.000000 94.200000 0.840000 ;
      RECT 91.640000 0.000000 92.820000 0.840000 ;
      RECT 90.260000 0.000000 90.980000 0.840000 ;
      RECT 88.880000 0.000000 89.600000 0.840000 ;
      RECT 87.040000 0.000000 88.220000 0.840000 ;
      RECT 85.660000 0.000000 86.380000 0.840000 ;
      RECT 84.280000 0.000000 85.000000 0.840000 ;
      RECT 82.900000 0.000000 83.620000 0.840000 ;
      RECT 81.060000 0.000000 82.240000 0.840000 ;
      RECT 79.680000 0.000000 80.400000 0.840000 ;
      RECT 78.300000 0.000000 79.020000 0.840000 ;
      RECT 76.460000 0.000000 77.640000 0.840000 ;
      RECT 75.080000 0.000000 75.800000 0.840000 ;
      RECT 73.700000 0.000000 74.420000 0.840000 ;
      RECT 72.320000 0.000000 73.040000 0.840000 ;
      RECT 70.480000 0.000000 71.660000 0.840000 ;
      RECT 69.100000 0.000000 69.820000 0.840000 ;
      RECT 67.720000 0.000000 68.440000 0.840000 ;
      RECT 65.880000 0.000000 67.060000 0.840000 ;
      RECT 64.500000 0.000000 65.220000 0.840000 ;
      RECT 63.120000 0.000000 63.840000 0.840000 ;
      RECT 61.280000 0.000000 62.460000 0.840000 ;
      RECT 59.900000 0.000000 60.620000 0.840000 ;
      RECT 58.520000 0.000000 59.240000 0.840000 ;
      RECT 57.140000 0.000000 57.860000 0.840000 ;
      RECT 55.300000 0.000000 56.480000 0.840000 ;
      RECT 53.920000 0.000000 54.640000 0.840000 ;
      RECT 52.540000 0.000000 53.260000 0.840000 ;
      RECT 50.700000 0.000000 51.880000 0.840000 ;
      RECT 49.320000 0.000000 50.040000 0.840000 ;
      RECT 47.940000 0.000000 48.660000 0.840000 ;
      RECT 46.100000 0.000000 47.280000 0.840000 ;
      RECT 44.720000 0.000000 45.440000 0.840000 ;
      RECT 43.340000 0.000000 44.060000 0.840000 ;
      RECT 41.960000 0.000000 42.680000 0.840000 ;
      RECT 40.120000 0.000000 41.300000 0.840000 ;
      RECT 38.740000 0.000000 39.460000 0.840000 ;
      RECT 37.360000 0.000000 38.080000 0.840000 ;
      RECT 35.520000 0.000000 36.700000 0.840000 ;
      RECT 34.140000 0.000000 34.860000 0.840000 ;
      RECT 32.760000 0.000000 33.480000 0.840000 ;
      RECT 31.380000 0.000000 32.100000 0.840000 ;
      RECT 29.540000 0.000000 30.720000 0.840000 ;
      RECT 28.160000 0.000000 28.880000 0.840000 ;
      RECT 26.780000 0.000000 27.500000 0.840000 ;
      RECT 24.940000 0.000000 26.120000 0.840000 ;
      RECT 23.560000 0.000000 24.280000 0.840000 ;
      RECT 22.180000 0.000000 22.900000 0.840000 ;
      RECT 20.340000 0.000000 21.520000 0.840000 ;
      RECT 18.960000 0.000000 19.680000 0.840000 ;
      RECT 17.580000 0.000000 18.300000 0.840000 ;
      RECT 16.200000 0.000000 16.920000 0.840000 ;
      RECT 14.360000 0.000000 15.540000 0.840000 ;
      RECT 12.980000 0.000000 13.700000 0.840000 ;
      RECT 11.600000 0.000000 12.320000 0.840000 ;
      RECT 9.760000 0.000000 10.940000 0.840000 ;
      RECT 8.380000 0.000000 9.100000 0.840000 ;
      RECT 7.000000 0.000000 7.720000 0.840000 ;
      RECT 5.620000 0.000000 6.340000 0.840000 ;
      RECT 0.000000 0.000000 4.960000 0.840000 ;
    LAYER met3 ;
      RECT 0.000000 198.320000 200.100000 200.260000 ;
      RECT 1.000000 193.880000 199.100000 194.720000 ;
      RECT 0.000000 193.320000 200.100000 193.880000 ;
      RECT 199.370000 193.030000 200.100000 193.320000 ;
      RECT 0.000000 193.030000 0.730000 193.320000 ;
      RECT 186.560000 192.240000 197.570000 193.320000 ;
      RECT 141.560000 192.240000 184.760000 193.320000 ;
      RECT 96.560000 192.240000 139.760000 193.320000 ;
      RECT 51.560000 192.240000 94.760000 193.320000 ;
      RECT 6.560000 192.240000 49.760000 193.320000 ;
      RECT 2.530000 192.240000 4.595000 193.320000 ;
      RECT 1.000000 192.050000 199.100000 192.240000 ;
      RECT 0.000000 191.810000 200.100000 192.050000 ;
      RECT 1.000000 190.830000 199.100000 191.810000 ;
      RECT 0.000000 190.600000 200.100000 190.830000 ;
      RECT 197.570000 189.980000 200.100000 190.600000 ;
      RECT 0.000000 189.980000 2.530000 190.600000 ;
      RECT 197.570000 189.520000 199.100000 189.980000 ;
      RECT 188.560000 189.520000 195.770000 190.600000 ;
      RECT 143.560000 189.520000 186.760000 190.600000 ;
      RECT 98.560000 189.520000 141.760000 190.600000 ;
      RECT 53.560000 189.520000 96.760000 190.600000 ;
      RECT 8.560000 189.520000 51.760000 190.600000 ;
      RECT 4.330000 189.520000 6.760000 190.600000 ;
      RECT 1.000000 189.520000 2.530000 189.980000 ;
      RECT 1.000000 189.000000 199.100000 189.520000 ;
      RECT 0.000000 188.760000 200.100000 189.000000 ;
      RECT 1.000000 187.880000 199.100000 188.760000 ;
      RECT 199.370000 186.930000 200.100000 187.780000 ;
      RECT 0.000000 186.930000 0.730000 187.780000 ;
      RECT 186.560000 186.800000 197.570000 187.880000 ;
      RECT 141.560000 186.800000 184.760000 187.880000 ;
      RECT 96.560000 186.800000 139.760000 187.880000 ;
      RECT 51.560000 186.800000 94.760000 187.880000 ;
      RECT 6.560000 186.800000 49.760000 187.880000 ;
      RECT 2.530000 186.800000 4.595000 187.880000 ;
      RECT 1.000000 185.950000 199.100000 186.800000 ;
      RECT 0.000000 185.710000 200.100000 185.950000 ;
      RECT 1.000000 185.160000 199.100000 185.710000 ;
      RECT 197.570000 184.730000 199.100000 185.160000 ;
      RECT 1.000000 184.730000 2.530000 185.160000 ;
      RECT 197.570000 184.080000 200.100000 184.730000 ;
      RECT 188.560000 184.080000 195.770000 185.160000 ;
      RECT 143.560000 184.080000 186.760000 185.160000 ;
      RECT 98.560000 184.080000 141.760000 185.160000 ;
      RECT 53.560000 184.080000 96.760000 185.160000 ;
      RECT 8.560000 184.080000 51.760000 185.160000 ;
      RECT 4.330000 184.080000 6.760000 185.160000 ;
      RECT 0.000000 184.080000 2.530000 184.730000 ;
      RECT 0.000000 183.880000 200.100000 184.080000 ;
      RECT 1.000000 182.900000 199.100000 183.880000 ;
      RECT 0.000000 182.660000 200.100000 182.900000 ;
      RECT 1.000000 182.440000 199.100000 182.660000 ;
      RECT 199.370000 181.440000 200.100000 181.680000 ;
      RECT 0.000000 181.440000 0.730000 181.680000 ;
      RECT 186.560000 181.360000 197.570000 182.440000 ;
      RECT 141.560000 181.360000 184.760000 182.440000 ;
      RECT 96.560000 181.360000 139.760000 182.440000 ;
      RECT 51.560000 181.360000 94.760000 182.440000 ;
      RECT 6.560000 181.360000 49.760000 182.440000 ;
      RECT 2.530000 181.360000 4.595000 182.440000 ;
      RECT 1.000000 180.460000 199.100000 181.360000 ;
      RECT 0.000000 179.720000 200.100000 180.460000 ;
      RECT 197.570000 179.610000 200.100000 179.720000 ;
      RECT 0.000000 179.610000 2.530000 179.720000 ;
      RECT 197.570000 178.640000 199.100000 179.610000 ;
      RECT 188.560000 178.640000 195.770000 179.720000 ;
      RECT 143.560000 178.640000 186.760000 179.720000 ;
      RECT 98.560000 178.640000 141.760000 179.720000 ;
      RECT 53.560000 178.640000 96.760000 179.720000 ;
      RECT 8.560000 178.640000 51.760000 179.720000 ;
      RECT 4.330000 178.640000 6.760000 179.720000 ;
      RECT 1.000000 178.640000 2.530000 179.610000 ;
      RECT 1.000000 178.630000 199.100000 178.640000 ;
      RECT 0.000000 178.390000 200.100000 178.630000 ;
      RECT 1.000000 177.410000 199.100000 178.390000 ;
      RECT 0.000000 177.000000 200.100000 177.410000 ;
      RECT 199.370000 176.560000 200.100000 177.000000 ;
      RECT 0.000000 176.560000 0.730000 177.000000 ;
      RECT 186.560000 175.920000 197.570000 177.000000 ;
      RECT 141.560000 175.920000 184.760000 177.000000 ;
      RECT 96.560000 175.920000 139.760000 177.000000 ;
      RECT 51.560000 175.920000 94.760000 177.000000 ;
      RECT 6.560000 175.920000 49.760000 177.000000 ;
      RECT 2.530000 175.920000 4.595000 177.000000 ;
      RECT 1.000000 175.580000 199.100000 175.920000 ;
      RECT 0.000000 175.340000 200.100000 175.580000 ;
      RECT 1.000000 174.360000 199.100000 175.340000 ;
      RECT 0.000000 174.280000 200.100000 174.360000 ;
      RECT 197.570000 173.510000 200.100000 174.280000 ;
      RECT 0.000000 173.510000 2.530000 174.280000 ;
      RECT 197.570000 173.200000 199.100000 173.510000 ;
      RECT 188.560000 173.200000 195.770000 174.280000 ;
      RECT 143.560000 173.200000 186.760000 174.280000 ;
      RECT 98.560000 173.200000 141.760000 174.280000 ;
      RECT 53.560000 173.200000 96.760000 174.280000 ;
      RECT 8.560000 173.200000 51.760000 174.280000 ;
      RECT 4.330000 173.200000 6.760000 174.280000 ;
      RECT 1.000000 173.200000 2.530000 173.510000 ;
      RECT 1.000000 172.530000 199.100000 173.200000 ;
      RECT 0.000000 172.290000 200.100000 172.530000 ;
      RECT 1.000000 171.560000 199.100000 172.290000 ;
      RECT 199.370000 170.480000 200.100000 171.310000 ;
      RECT 186.560000 170.480000 197.570000 171.560000 ;
      RECT 141.560000 170.480000 184.760000 171.560000 ;
      RECT 96.560000 170.480000 139.760000 171.560000 ;
      RECT 51.560000 170.480000 94.760000 171.560000 ;
      RECT 6.560000 170.480000 49.760000 171.560000 ;
      RECT 2.530000 170.480000 4.595000 171.560000 ;
      RECT 0.000000 170.480000 0.730000 171.310000 ;
      RECT 0.000000 170.460000 200.100000 170.480000 ;
      RECT 1.000000 169.480000 199.100000 170.460000 ;
      RECT 0.000000 169.240000 200.100000 169.480000 ;
      RECT 1.000000 168.840000 199.100000 169.240000 ;
      RECT 197.570000 168.260000 199.100000 168.840000 ;
      RECT 1.000000 168.260000 2.530000 168.840000 ;
      RECT 197.570000 168.020000 200.100000 168.260000 ;
      RECT 0.000000 168.020000 2.530000 168.260000 ;
      RECT 197.570000 167.760000 199.100000 168.020000 ;
      RECT 188.560000 167.760000 195.770000 168.840000 ;
      RECT 143.560000 167.760000 186.760000 168.840000 ;
      RECT 98.560000 167.760000 141.760000 168.840000 ;
      RECT 53.560000 167.760000 96.760000 168.840000 ;
      RECT 8.560000 167.760000 51.760000 168.840000 ;
      RECT 4.330000 167.760000 6.760000 168.840000 ;
      RECT 1.000000 167.760000 2.530000 168.020000 ;
      RECT 1.000000 167.040000 199.100000 167.760000 ;
      RECT 0.000000 166.190000 200.100000 167.040000 ;
      RECT 1.000000 166.120000 199.100000 166.190000 ;
      RECT 199.370000 165.040000 200.100000 165.210000 ;
      RECT 186.560000 165.040000 197.570000 166.120000 ;
      RECT 141.560000 165.040000 184.760000 166.120000 ;
      RECT 96.560000 165.040000 139.760000 166.120000 ;
      RECT 51.560000 165.040000 94.760000 166.120000 ;
      RECT 6.560000 165.040000 49.760000 166.120000 ;
      RECT 2.530000 165.040000 4.595000 166.120000 ;
      RECT 0.000000 165.040000 0.730000 165.210000 ;
      RECT 0.000000 164.970000 200.100000 165.040000 ;
      RECT 1.000000 163.990000 199.100000 164.970000 ;
      RECT 0.000000 163.400000 200.100000 163.990000 ;
      RECT 197.570000 163.140000 200.100000 163.400000 ;
      RECT 0.000000 163.140000 2.530000 163.400000 ;
      RECT 197.570000 162.320000 199.100000 163.140000 ;
      RECT 188.560000 162.320000 195.770000 163.400000 ;
      RECT 143.560000 162.320000 186.760000 163.400000 ;
      RECT 98.560000 162.320000 141.760000 163.400000 ;
      RECT 53.560000 162.320000 96.760000 163.400000 ;
      RECT 8.560000 162.320000 51.760000 163.400000 ;
      RECT 4.330000 162.320000 6.760000 163.400000 ;
      RECT 1.000000 162.320000 2.530000 163.140000 ;
      RECT 1.000000 162.160000 199.100000 162.320000 ;
      RECT 0.000000 161.920000 200.100000 162.160000 ;
      RECT 1.000000 160.940000 199.100000 161.920000 ;
      RECT 0.000000 160.680000 200.100000 160.940000 ;
      RECT 199.370000 160.090000 200.100000 160.680000 ;
      RECT 0.000000 160.090000 0.730000 160.680000 ;
      RECT 186.560000 159.600000 197.570000 160.680000 ;
      RECT 141.560000 159.600000 184.760000 160.680000 ;
      RECT 96.560000 159.600000 139.760000 160.680000 ;
      RECT 51.560000 159.600000 94.760000 160.680000 ;
      RECT 6.560000 159.600000 49.760000 160.680000 ;
      RECT 2.530000 159.600000 4.595000 160.680000 ;
      RECT 1.000000 159.110000 199.100000 159.600000 ;
      RECT 0.000000 158.870000 200.100000 159.110000 ;
      RECT 1.000000 157.960000 199.100000 158.870000 ;
      RECT 197.570000 157.890000 199.100000 157.960000 ;
      RECT 1.000000 157.890000 2.530000 157.960000 ;
      RECT 197.570000 157.040000 200.100000 157.890000 ;
      RECT 0.000000 157.040000 2.530000 157.890000 ;
      RECT 197.570000 156.880000 199.100000 157.040000 ;
      RECT 188.560000 156.880000 195.770000 157.960000 ;
      RECT 143.560000 156.880000 186.760000 157.960000 ;
      RECT 98.560000 156.880000 141.760000 157.960000 ;
      RECT 53.560000 156.880000 96.760000 157.960000 ;
      RECT 8.560000 156.880000 51.760000 157.960000 ;
      RECT 4.330000 156.880000 6.760000 157.960000 ;
      RECT 1.000000 156.880000 2.530000 157.040000 ;
      RECT 1.000000 156.060000 199.100000 156.880000 ;
      RECT 0.000000 155.820000 200.100000 156.060000 ;
      RECT 1.000000 155.240000 199.100000 155.820000 ;
      RECT 199.370000 154.600000 200.100000 154.840000 ;
      RECT 0.000000 154.600000 0.730000 154.840000 ;
      RECT 186.560000 154.160000 197.570000 155.240000 ;
      RECT 141.560000 154.160000 184.760000 155.240000 ;
      RECT 96.560000 154.160000 139.760000 155.240000 ;
      RECT 51.560000 154.160000 94.760000 155.240000 ;
      RECT 6.560000 154.160000 49.760000 155.240000 ;
      RECT 2.530000 154.160000 4.595000 155.240000 ;
      RECT 1.000000 153.620000 199.100000 154.160000 ;
      RECT 0.000000 152.770000 200.100000 153.620000 ;
      RECT 1.000000 152.520000 199.100000 152.770000 ;
      RECT 197.570000 151.790000 199.100000 152.520000 ;
      RECT 1.000000 151.790000 2.530000 152.520000 ;
      RECT 197.570000 151.550000 200.100000 151.790000 ;
      RECT 0.000000 151.550000 2.530000 151.790000 ;
      RECT 197.570000 151.440000 199.100000 151.550000 ;
      RECT 188.560000 151.440000 195.770000 152.520000 ;
      RECT 143.560000 151.440000 186.760000 152.520000 ;
      RECT 98.560000 151.440000 141.760000 152.520000 ;
      RECT 53.560000 151.440000 96.760000 152.520000 ;
      RECT 8.560000 151.440000 51.760000 152.520000 ;
      RECT 4.330000 151.440000 6.760000 152.520000 ;
      RECT 1.000000 151.440000 2.530000 151.550000 ;
      RECT 1.000000 150.570000 199.100000 151.440000 ;
      RECT 0.000000 149.800000 200.100000 150.570000 ;
      RECT 199.370000 149.720000 200.100000 149.800000 ;
      RECT 0.000000 149.720000 0.730000 149.800000 ;
      RECT 199.370000 148.720000 200.100000 148.740000 ;
      RECT 186.560000 148.720000 197.570000 149.800000 ;
      RECT 141.560000 148.720000 184.760000 149.800000 ;
      RECT 96.560000 148.720000 139.760000 149.800000 ;
      RECT 51.560000 148.720000 94.760000 149.800000 ;
      RECT 6.560000 148.720000 49.760000 149.800000 ;
      RECT 2.530000 148.720000 4.595000 149.800000 ;
      RECT 0.000000 148.720000 0.730000 148.740000 ;
      RECT 0.000000 148.500000 200.100000 148.720000 ;
      RECT 1.000000 147.520000 199.100000 148.500000 ;
      RECT 0.000000 147.080000 200.100000 147.520000 ;
      RECT 197.570000 146.670000 200.100000 147.080000 ;
      RECT 0.000000 146.670000 2.530000 147.080000 ;
      RECT 197.570000 146.000000 199.100000 146.670000 ;
      RECT 188.560000 146.000000 195.770000 147.080000 ;
      RECT 143.560000 146.000000 186.760000 147.080000 ;
      RECT 98.560000 146.000000 141.760000 147.080000 ;
      RECT 53.560000 146.000000 96.760000 147.080000 ;
      RECT 8.560000 146.000000 51.760000 147.080000 ;
      RECT 4.330000 146.000000 6.760000 147.080000 ;
      RECT 1.000000 146.000000 2.530000 146.670000 ;
      RECT 1.000000 145.690000 199.100000 146.000000 ;
      RECT 0.000000 145.450000 200.100000 145.690000 ;
      RECT 1.000000 144.470000 199.100000 145.450000 ;
      RECT 0.000000 144.360000 200.100000 144.470000 ;
      RECT 199.370000 144.230000 200.100000 144.360000 ;
      RECT 0.000000 144.230000 0.730000 144.360000 ;
      RECT 186.560000 143.280000 197.570000 144.360000 ;
      RECT 141.560000 143.280000 184.760000 144.360000 ;
      RECT 96.560000 143.280000 139.760000 144.360000 ;
      RECT 51.560000 143.280000 94.760000 144.360000 ;
      RECT 6.560000 143.280000 49.760000 144.360000 ;
      RECT 2.530000 143.280000 4.595000 144.360000 ;
      RECT 1.000000 143.250000 199.100000 143.280000 ;
      RECT 0.000000 142.400000 200.100000 143.250000 ;
      RECT 1.000000 141.640000 199.100000 142.400000 ;
      RECT 197.570000 141.420000 199.100000 141.640000 ;
      RECT 1.000000 141.420000 2.530000 141.640000 ;
      RECT 197.570000 141.180000 200.100000 141.420000 ;
      RECT 0.000000 141.180000 2.530000 141.420000 ;
      RECT 197.570000 140.560000 199.100000 141.180000 ;
      RECT 188.560000 140.560000 195.770000 141.640000 ;
      RECT 143.560000 140.560000 186.760000 141.640000 ;
      RECT 98.560000 140.560000 141.760000 141.640000 ;
      RECT 53.560000 140.560000 96.760000 141.640000 ;
      RECT 8.560000 140.560000 51.760000 141.640000 ;
      RECT 4.330000 140.560000 6.760000 141.640000 ;
      RECT 1.000000 140.560000 2.530000 141.180000 ;
      RECT 1.000000 140.200000 199.100000 140.560000 ;
      RECT 0.000000 139.350000 200.100000 140.200000 ;
      RECT 1.000000 138.920000 199.100000 139.350000 ;
      RECT 199.370000 138.130000 200.100000 138.370000 ;
      RECT 0.000000 138.130000 0.730000 138.370000 ;
      RECT 186.560000 137.840000 197.570000 138.920000 ;
      RECT 141.560000 137.840000 184.760000 138.920000 ;
      RECT 96.560000 137.840000 139.760000 138.920000 ;
      RECT 51.560000 137.840000 94.760000 138.920000 ;
      RECT 6.560000 137.840000 49.760000 138.920000 ;
      RECT 2.530000 137.840000 4.595000 138.920000 ;
      RECT 1.000000 137.150000 199.100000 137.840000 ;
      RECT 0.000000 136.300000 200.100000 137.150000 ;
      RECT 1.000000 136.200000 199.100000 136.300000 ;
      RECT 197.570000 135.320000 199.100000 136.200000 ;
      RECT 1.000000 135.320000 2.530000 136.200000 ;
      RECT 197.570000 135.120000 200.100000 135.320000 ;
      RECT 188.560000 135.120000 195.770000 136.200000 ;
      RECT 143.560000 135.120000 186.760000 136.200000 ;
      RECT 98.560000 135.120000 141.760000 136.200000 ;
      RECT 53.560000 135.120000 96.760000 136.200000 ;
      RECT 8.560000 135.120000 51.760000 136.200000 ;
      RECT 4.330000 135.120000 6.760000 136.200000 ;
      RECT 0.000000 135.120000 2.530000 135.320000 ;
      RECT 0.000000 135.080000 200.100000 135.120000 ;
      RECT 1.000000 134.100000 199.100000 135.080000 ;
      RECT 0.000000 133.480000 200.100000 134.100000 ;
      RECT 199.370000 133.250000 200.100000 133.480000 ;
      RECT 0.000000 133.250000 0.730000 133.480000 ;
      RECT 186.560000 132.400000 197.570000 133.480000 ;
      RECT 141.560000 132.400000 184.760000 133.480000 ;
      RECT 96.560000 132.400000 139.760000 133.480000 ;
      RECT 51.560000 132.400000 94.760000 133.480000 ;
      RECT 6.560000 132.400000 49.760000 133.480000 ;
      RECT 2.530000 132.400000 4.595000 133.480000 ;
      RECT 1.000000 132.270000 199.100000 132.400000 ;
      RECT 0.000000 132.030000 200.100000 132.270000 ;
      RECT 1.000000 131.050000 199.100000 132.030000 ;
      RECT 0.000000 130.810000 200.100000 131.050000 ;
      RECT 1.000000 130.760000 199.100000 130.810000 ;
      RECT 197.570000 129.830000 199.100000 130.760000 ;
      RECT 1.000000 129.830000 2.530000 130.760000 ;
      RECT 197.570000 129.680000 200.100000 129.830000 ;
      RECT 188.560000 129.680000 195.770000 130.760000 ;
      RECT 143.560000 129.680000 186.760000 130.760000 ;
      RECT 98.560000 129.680000 141.760000 130.760000 ;
      RECT 53.560000 129.680000 96.760000 130.760000 ;
      RECT 8.560000 129.680000 51.760000 130.760000 ;
      RECT 4.330000 129.680000 6.760000 130.760000 ;
      RECT 0.000000 129.680000 2.530000 129.830000 ;
      RECT 0.000000 128.980000 200.100000 129.680000 ;
      RECT 1.000000 128.040000 199.100000 128.980000 ;
      RECT 199.370000 127.760000 200.100000 128.000000 ;
      RECT 0.000000 127.760000 0.730000 128.000000 ;
      RECT 186.560000 126.960000 197.570000 128.040000 ;
      RECT 141.560000 126.960000 184.760000 128.040000 ;
      RECT 96.560000 126.960000 139.760000 128.040000 ;
      RECT 51.560000 126.960000 94.760000 128.040000 ;
      RECT 6.560000 126.960000 49.760000 128.040000 ;
      RECT 2.530000 126.960000 4.595000 128.040000 ;
      RECT 1.000000 126.780000 199.100000 126.960000 ;
      RECT 0.000000 125.930000 200.100000 126.780000 ;
      RECT 1.000000 125.320000 199.100000 125.930000 ;
      RECT 197.570000 124.950000 199.100000 125.320000 ;
      RECT 1.000000 124.950000 2.530000 125.320000 ;
      RECT 197.570000 124.710000 200.100000 124.950000 ;
      RECT 0.000000 124.710000 2.530000 124.950000 ;
      RECT 197.570000 124.240000 199.100000 124.710000 ;
      RECT 188.560000 124.240000 195.770000 125.320000 ;
      RECT 143.560000 124.240000 186.760000 125.320000 ;
      RECT 98.560000 124.240000 141.760000 125.320000 ;
      RECT 53.560000 124.240000 96.760000 125.320000 ;
      RECT 8.560000 124.240000 51.760000 125.320000 ;
      RECT 4.330000 124.240000 6.760000 125.320000 ;
      RECT 1.000000 124.240000 2.530000 124.710000 ;
      RECT 1.000000 123.730000 199.100000 124.240000 ;
      RECT 0.000000 122.880000 200.100000 123.730000 ;
      RECT 1.000000 122.600000 199.100000 122.880000 ;
      RECT 199.370000 121.660000 200.100000 121.900000 ;
      RECT 0.000000 121.660000 0.730000 121.900000 ;
      RECT 186.560000 121.520000 197.570000 122.600000 ;
      RECT 141.560000 121.520000 184.760000 122.600000 ;
      RECT 96.560000 121.520000 139.760000 122.600000 ;
      RECT 51.560000 121.520000 94.760000 122.600000 ;
      RECT 6.560000 121.520000 49.760000 122.600000 ;
      RECT 2.530000 121.520000 4.595000 122.600000 ;
      RECT 1.000000 120.680000 199.100000 121.520000 ;
      RECT 0.000000 119.880000 200.100000 120.680000 ;
      RECT 197.570000 119.830000 200.100000 119.880000 ;
      RECT 0.000000 119.830000 2.530000 119.880000 ;
      RECT 197.570000 118.850000 199.100000 119.830000 ;
      RECT 1.000000 118.850000 2.530000 119.830000 ;
      RECT 197.570000 118.800000 200.100000 118.850000 ;
      RECT 188.560000 118.800000 195.770000 119.880000 ;
      RECT 143.560000 118.800000 186.760000 119.880000 ;
      RECT 98.560000 118.800000 141.760000 119.880000 ;
      RECT 53.560000 118.800000 96.760000 119.880000 ;
      RECT 8.560000 118.800000 51.760000 119.880000 ;
      RECT 4.330000 118.800000 6.760000 119.880000 ;
      RECT 0.000000 118.800000 2.530000 118.850000 ;
      RECT 0.000000 118.610000 200.100000 118.800000 ;
      RECT 1.000000 117.630000 199.100000 118.610000 ;
      RECT 0.000000 117.390000 200.100000 117.630000 ;
      RECT 1.000000 117.160000 199.100000 117.390000 ;
      RECT 199.370000 116.080000 200.100000 116.410000 ;
      RECT 186.560000 116.080000 197.570000 117.160000 ;
      RECT 141.560000 116.080000 184.760000 117.160000 ;
      RECT 96.560000 116.080000 139.760000 117.160000 ;
      RECT 51.560000 116.080000 94.760000 117.160000 ;
      RECT 6.560000 116.080000 49.760000 117.160000 ;
      RECT 2.530000 116.080000 4.595000 117.160000 ;
      RECT 0.000000 116.080000 0.730000 116.410000 ;
      RECT 0.000000 115.560000 200.100000 116.080000 ;
      RECT 1.000000 114.580000 199.100000 115.560000 ;
      RECT 0.000000 114.440000 200.100000 114.580000 ;
      RECT 197.570000 114.340000 200.100000 114.440000 ;
      RECT 0.000000 114.340000 2.530000 114.440000 ;
      RECT 197.570000 113.360000 199.100000 114.340000 ;
      RECT 188.560000 113.360000 195.770000 114.440000 ;
      RECT 143.560000 113.360000 186.760000 114.440000 ;
      RECT 98.560000 113.360000 141.760000 114.440000 ;
      RECT 53.560000 113.360000 96.760000 114.440000 ;
      RECT 8.560000 113.360000 51.760000 114.440000 ;
      RECT 4.330000 113.360000 6.760000 114.440000 ;
      RECT 1.000000 113.360000 2.530000 114.340000 ;
      RECT 0.000000 112.510000 200.100000 113.360000 ;
      RECT 1.000000 111.720000 199.100000 112.510000 ;
      RECT 199.370000 111.290000 200.100000 111.530000 ;
      RECT 0.000000 111.290000 0.730000 111.530000 ;
      RECT 186.560000 110.640000 197.570000 111.720000 ;
      RECT 141.560000 110.640000 184.760000 111.720000 ;
      RECT 96.560000 110.640000 139.760000 111.720000 ;
      RECT 51.560000 110.640000 94.760000 111.720000 ;
      RECT 6.560000 110.640000 49.760000 111.720000 ;
      RECT 2.530000 110.640000 4.595000 111.720000 ;
      RECT 1.000000 110.310000 199.100000 110.640000 ;
      RECT 0.000000 109.460000 200.100000 110.310000 ;
      RECT 1.000000 109.000000 199.100000 109.460000 ;
      RECT 197.570000 108.480000 199.100000 109.000000 ;
      RECT 1.000000 108.480000 2.530000 109.000000 ;
      RECT 197.570000 108.240000 200.100000 108.480000 ;
      RECT 0.000000 108.240000 2.530000 108.480000 ;
      RECT 197.570000 107.920000 199.100000 108.240000 ;
      RECT 188.560000 107.920000 195.770000 109.000000 ;
      RECT 143.560000 107.920000 186.760000 109.000000 ;
      RECT 98.560000 107.920000 141.760000 109.000000 ;
      RECT 53.560000 107.920000 96.760000 109.000000 ;
      RECT 8.560000 107.920000 51.760000 109.000000 ;
      RECT 4.330000 107.920000 6.760000 109.000000 ;
      RECT 1.000000 107.920000 2.530000 108.240000 ;
      RECT 1.000000 107.260000 199.100000 107.920000 ;
      RECT 0.000000 106.410000 200.100000 107.260000 ;
      RECT 1.000000 106.280000 199.100000 106.410000 ;
      RECT 199.370000 105.200000 200.100000 105.430000 ;
      RECT 186.560000 105.200000 197.570000 106.280000 ;
      RECT 141.560000 105.200000 184.760000 106.280000 ;
      RECT 96.560000 105.200000 139.760000 106.280000 ;
      RECT 51.560000 105.200000 94.760000 106.280000 ;
      RECT 6.560000 105.200000 49.760000 106.280000 ;
      RECT 2.530000 105.200000 4.595000 106.280000 ;
      RECT 0.000000 105.200000 0.730000 105.430000 ;
      RECT 0.000000 105.190000 200.100000 105.200000 ;
      RECT 1.000000 104.210000 199.100000 105.190000 ;
      RECT 0.000000 103.970000 200.100000 104.210000 ;
      RECT 1.000000 103.560000 199.100000 103.970000 ;
      RECT 197.570000 102.990000 199.100000 103.560000 ;
      RECT 1.000000 102.990000 2.530000 103.560000 ;
      RECT 197.570000 102.480000 200.100000 102.990000 ;
      RECT 188.560000 102.480000 195.770000 103.560000 ;
      RECT 143.560000 102.480000 186.760000 103.560000 ;
      RECT 98.560000 102.480000 141.760000 103.560000 ;
      RECT 53.560000 102.480000 96.760000 103.560000 ;
      RECT 8.560000 102.480000 51.760000 103.560000 ;
      RECT 4.330000 102.480000 6.760000 103.560000 ;
      RECT 0.000000 102.480000 2.530000 102.990000 ;
      RECT 0.000000 102.140000 200.100000 102.480000 ;
      RECT 1.000000 101.160000 199.100000 102.140000 ;
      RECT 0.000000 100.920000 200.100000 101.160000 ;
      RECT 1.000000 100.840000 199.100000 100.920000 ;
      RECT 199.370000 99.760000 200.100000 99.940000 ;
      RECT 186.560000 99.760000 197.570000 100.840000 ;
      RECT 141.560000 99.760000 184.760000 100.840000 ;
      RECT 96.560000 99.760000 139.760000 100.840000 ;
      RECT 51.560000 99.760000 94.760000 100.840000 ;
      RECT 6.560000 99.760000 49.760000 100.840000 ;
      RECT 2.530000 99.760000 4.595000 100.840000 ;
      RECT 0.000000 99.760000 0.730000 99.940000 ;
      RECT 0.000000 99.090000 200.100000 99.760000 ;
      RECT 1.000000 98.120000 199.100000 99.090000 ;
      RECT 197.570000 98.110000 199.100000 98.120000 ;
      RECT 1.000000 98.110000 2.530000 98.120000 ;
      RECT 197.570000 97.870000 200.100000 98.110000 ;
      RECT 0.000000 97.870000 2.530000 98.110000 ;
      RECT 197.570000 97.040000 199.100000 97.870000 ;
      RECT 188.560000 97.040000 195.770000 98.120000 ;
      RECT 143.560000 97.040000 186.760000 98.120000 ;
      RECT 98.560000 97.040000 141.760000 98.120000 ;
      RECT 53.560000 97.040000 96.760000 98.120000 ;
      RECT 8.560000 97.040000 51.760000 98.120000 ;
      RECT 4.330000 97.040000 6.760000 98.120000 ;
      RECT 1.000000 97.040000 2.530000 97.870000 ;
      RECT 1.000000 96.890000 199.100000 97.040000 ;
      RECT 0.000000 96.040000 200.100000 96.890000 ;
      RECT 1.000000 95.400000 199.100000 96.040000 ;
      RECT 199.370000 94.820000 200.100000 95.060000 ;
      RECT 0.000000 94.820000 0.730000 95.060000 ;
      RECT 186.560000 94.320000 197.570000 95.400000 ;
      RECT 141.560000 94.320000 184.760000 95.400000 ;
      RECT 96.560000 94.320000 139.760000 95.400000 ;
      RECT 51.560000 94.320000 94.760000 95.400000 ;
      RECT 6.560000 94.320000 49.760000 95.400000 ;
      RECT 2.530000 94.320000 4.595000 95.400000 ;
      RECT 1.000000 93.840000 199.100000 94.320000 ;
      RECT 0.000000 93.600000 200.100000 93.840000 ;
      RECT 1.000000 92.680000 199.100000 93.600000 ;
      RECT 197.570000 92.620000 199.100000 92.680000 ;
      RECT 1.000000 92.620000 2.530000 92.680000 ;
      RECT 197.570000 91.770000 200.100000 92.620000 ;
      RECT 0.000000 91.770000 2.530000 92.620000 ;
      RECT 197.570000 91.600000 199.100000 91.770000 ;
      RECT 188.560000 91.600000 195.770000 92.680000 ;
      RECT 143.560000 91.600000 186.760000 92.680000 ;
      RECT 98.560000 91.600000 141.760000 92.680000 ;
      RECT 53.560000 91.600000 96.760000 92.680000 ;
      RECT 8.560000 91.600000 51.760000 92.680000 ;
      RECT 4.330000 91.600000 6.760000 92.680000 ;
      RECT 1.000000 91.600000 2.530000 91.770000 ;
      RECT 1.000000 90.790000 199.100000 91.600000 ;
      RECT 0.000000 90.550000 200.100000 90.790000 ;
      RECT 1.000000 89.960000 199.100000 90.550000 ;
      RECT 199.370000 88.880000 200.100000 89.570000 ;
      RECT 186.560000 88.880000 197.570000 89.960000 ;
      RECT 141.560000 88.880000 184.760000 89.960000 ;
      RECT 96.560000 88.880000 139.760000 89.960000 ;
      RECT 51.560000 88.880000 94.760000 89.960000 ;
      RECT 6.560000 88.880000 49.760000 89.960000 ;
      RECT 2.530000 88.880000 4.595000 89.960000 ;
      RECT 0.000000 88.880000 0.730000 89.570000 ;
      RECT 0.000000 88.720000 200.100000 88.880000 ;
      RECT 1.000000 87.740000 199.100000 88.720000 ;
      RECT 0.000000 87.500000 200.100000 87.740000 ;
      RECT 1.000000 87.240000 199.100000 87.500000 ;
      RECT 197.570000 86.520000 199.100000 87.240000 ;
      RECT 1.000000 86.520000 2.530000 87.240000 ;
      RECT 197.570000 86.160000 200.100000 86.520000 ;
      RECT 188.560000 86.160000 195.770000 87.240000 ;
      RECT 143.560000 86.160000 186.760000 87.240000 ;
      RECT 98.560000 86.160000 141.760000 87.240000 ;
      RECT 53.560000 86.160000 96.760000 87.240000 ;
      RECT 8.560000 86.160000 51.760000 87.240000 ;
      RECT 4.330000 86.160000 6.760000 87.240000 ;
      RECT 0.000000 86.160000 2.530000 86.520000 ;
      RECT 0.000000 85.670000 200.100000 86.160000 ;
      RECT 1.000000 84.690000 199.100000 85.670000 ;
      RECT 0.000000 84.520000 200.100000 84.690000 ;
      RECT 199.370000 84.450000 200.100000 84.520000 ;
      RECT 0.000000 84.450000 0.730000 84.520000 ;
      RECT 199.370000 83.440000 200.100000 83.470000 ;
      RECT 186.560000 83.440000 197.570000 84.520000 ;
      RECT 141.560000 83.440000 184.760000 84.520000 ;
      RECT 96.560000 83.440000 139.760000 84.520000 ;
      RECT 51.560000 83.440000 94.760000 84.520000 ;
      RECT 6.560000 83.440000 49.760000 84.520000 ;
      RECT 2.530000 83.440000 4.595000 84.520000 ;
      RECT 0.000000 83.440000 0.730000 83.470000 ;
      RECT 0.000000 82.620000 200.100000 83.440000 ;
      RECT 1.000000 81.800000 199.100000 82.620000 ;
      RECT 197.570000 81.640000 199.100000 81.800000 ;
      RECT 1.000000 81.640000 2.530000 81.800000 ;
      RECT 197.570000 81.400000 200.100000 81.640000 ;
      RECT 0.000000 81.400000 2.530000 81.640000 ;
      RECT 197.570000 80.720000 199.100000 81.400000 ;
      RECT 188.560000 80.720000 195.770000 81.800000 ;
      RECT 143.560000 80.720000 186.760000 81.800000 ;
      RECT 98.560000 80.720000 141.760000 81.800000 ;
      RECT 53.560000 80.720000 96.760000 81.800000 ;
      RECT 8.560000 80.720000 51.760000 81.800000 ;
      RECT 4.330000 80.720000 6.760000 81.800000 ;
      RECT 1.000000 80.720000 2.530000 81.400000 ;
      RECT 1.000000 80.420000 199.100000 80.720000 ;
      RECT 0.000000 80.180000 200.100000 80.420000 ;
      RECT 1.000000 79.200000 199.100000 80.180000 ;
      RECT 0.000000 79.080000 200.100000 79.200000 ;
      RECT 199.370000 78.350000 200.100000 79.080000 ;
      RECT 0.000000 78.350000 0.730000 79.080000 ;
      RECT 186.560000 78.000000 197.570000 79.080000 ;
      RECT 141.560000 78.000000 184.760000 79.080000 ;
      RECT 96.560000 78.000000 139.760000 79.080000 ;
      RECT 51.560000 78.000000 94.760000 79.080000 ;
      RECT 6.560000 78.000000 49.760000 79.080000 ;
      RECT 2.530000 78.000000 4.595000 79.080000 ;
      RECT 1.000000 77.370000 199.100000 78.000000 ;
      RECT 0.000000 77.130000 200.100000 77.370000 ;
      RECT 1.000000 76.360000 199.100000 77.130000 ;
      RECT 197.570000 76.150000 199.100000 76.360000 ;
      RECT 1.000000 76.150000 2.530000 76.360000 ;
      RECT 197.570000 75.300000 200.100000 76.150000 ;
      RECT 0.000000 75.300000 2.530000 76.150000 ;
      RECT 197.570000 75.280000 199.100000 75.300000 ;
      RECT 188.560000 75.280000 195.770000 76.360000 ;
      RECT 143.560000 75.280000 186.760000 76.360000 ;
      RECT 98.560000 75.280000 141.760000 76.360000 ;
      RECT 53.560000 75.280000 96.760000 76.360000 ;
      RECT 8.560000 75.280000 51.760000 76.360000 ;
      RECT 4.330000 75.280000 6.760000 76.360000 ;
      RECT 1.000000 75.280000 2.530000 75.300000 ;
      RECT 1.000000 74.320000 199.100000 75.280000 ;
      RECT 0.000000 74.080000 200.100000 74.320000 ;
      RECT 1.000000 73.640000 199.100000 74.080000 ;
      RECT 199.370000 72.560000 200.100000 73.100000 ;
      RECT 186.560000 72.560000 197.570000 73.640000 ;
      RECT 141.560000 72.560000 184.760000 73.640000 ;
      RECT 96.560000 72.560000 139.760000 73.640000 ;
      RECT 51.560000 72.560000 94.760000 73.640000 ;
      RECT 6.560000 72.560000 49.760000 73.640000 ;
      RECT 2.530000 72.560000 4.595000 73.640000 ;
      RECT 0.000000 72.560000 0.730000 73.100000 ;
      RECT 0.000000 72.250000 200.100000 72.560000 ;
      RECT 1.000000 71.270000 199.100000 72.250000 ;
      RECT 0.000000 71.030000 200.100000 71.270000 ;
      RECT 1.000000 70.920000 199.100000 71.030000 ;
      RECT 197.570000 70.050000 199.100000 70.920000 ;
      RECT 1.000000 70.050000 2.530000 70.920000 ;
      RECT 197.570000 69.840000 200.100000 70.050000 ;
      RECT 188.560000 69.840000 195.770000 70.920000 ;
      RECT 143.560000 69.840000 186.760000 70.920000 ;
      RECT 98.560000 69.840000 141.760000 70.920000 ;
      RECT 53.560000 69.840000 96.760000 70.920000 ;
      RECT 8.560000 69.840000 51.760000 70.920000 ;
      RECT 4.330000 69.840000 6.760000 70.920000 ;
      RECT 0.000000 69.840000 2.530000 70.050000 ;
      RECT 0.000000 69.200000 200.100000 69.840000 ;
      RECT 1.000000 68.220000 199.100000 69.200000 ;
      RECT 0.000000 68.200000 200.100000 68.220000 ;
      RECT 199.370000 67.980000 200.100000 68.200000 ;
      RECT 0.000000 67.980000 0.730000 68.200000 ;
      RECT 186.560000 67.120000 197.570000 68.200000 ;
      RECT 141.560000 67.120000 184.760000 68.200000 ;
      RECT 96.560000 67.120000 139.760000 68.200000 ;
      RECT 51.560000 67.120000 94.760000 68.200000 ;
      RECT 6.560000 67.120000 49.760000 68.200000 ;
      RECT 2.530000 67.120000 4.595000 68.200000 ;
      RECT 1.000000 67.000000 199.100000 67.120000 ;
      RECT 0.000000 66.760000 200.100000 67.000000 ;
      RECT 1.000000 65.780000 199.100000 66.760000 ;
      RECT 0.000000 65.480000 200.100000 65.780000 ;
      RECT 197.570000 64.930000 200.100000 65.480000 ;
      RECT 0.000000 64.930000 2.530000 65.480000 ;
      RECT 197.570000 64.400000 199.100000 64.930000 ;
      RECT 188.560000 64.400000 195.770000 65.480000 ;
      RECT 143.560000 64.400000 186.760000 65.480000 ;
      RECT 98.560000 64.400000 141.760000 65.480000 ;
      RECT 53.560000 64.400000 96.760000 65.480000 ;
      RECT 8.560000 64.400000 51.760000 65.480000 ;
      RECT 4.330000 64.400000 6.760000 65.480000 ;
      RECT 1.000000 64.400000 2.530000 64.930000 ;
      RECT 1.000000 63.950000 199.100000 64.400000 ;
      RECT 0.000000 63.710000 200.100000 63.950000 ;
      RECT 1.000000 62.760000 199.100000 63.710000 ;
      RECT 199.370000 61.880000 200.100000 62.730000 ;
      RECT 0.000000 61.880000 0.730000 62.730000 ;
      RECT 186.560000 61.680000 197.570000 62.760000 ;
      RECT 141.560000 61.680000 184.760000 62.760000 ;
      RECT 96.560000 61.680000 139.760000 62.760000 ;
      RECT 51.560000 61.680000 94.760000 62.760000 ;
      RECT 6.560000 61.680000 49.760000 62.760000 ;
      RECT 2.530000 61.680000 4.595000 62.760000 ;
      RECT 1.000000 60.900000 199.100000 61.680000 ;
      RECT 0.000000 60.660000 200.100000 60.900000 ;
      RECT 1.000000 60.040000 199.100000 60.660000 ;
      RECT 197.570000 59.680000 199.100000 60.040000 ;
      RECT 1.000000 59.680000 2.530000 60.040000 ;
      RECT 197.570000 58.960000 200.100000 59.680000 ;
      RECT 188.560000 58.960000 195.770000 60.040000 ;
      RECT 143.560000 58.960000 186.760000 60.040000 ;
      RECT 98.560000 58.960000 141.760000 60.040000 ;
      RECT 53.560000 58.960000 96.760000 60.040000 ;
      RECT 8.560000 58.960000 51.760000 60.040000 ;
      RECT 4.330000 58.960000 6.760000 60.040000 ;
      RECT 0.000000 58.960000 2.530000 59.680000 ;
      RECT 0.000000 58.830000 200.100000 58.960000 ;
      RECT 1.000000 57.850000 199.100000 58.830000 ;
      RECT 0.000000 57.610000 200.100000 57.850000 ;
      RECT 1.000000 57.320000 199.100000 57.610000 ;
      RECT 199.370000 56.240000 200.100000 56.630000 ;
      RECT 186.560000 56.240000 197.570000 57.320000 ;
      RECT 141.560000 56.240000 184.760000 57.320000 ;
      RECT 96.560000 56.240000 139.760000 57.320000 ;
      RECT 51.560000 56.240000 94.760000 57.320000 ;
      RECT 6.560000 56.240000 49.760000 57.320000 ;
      RECT 2.530000 56.240000 4.595000 57.320000 ;
      RECT 0.000000 56.240000 0.730000 56.630000 ;
      RECT 0.000000 55.780000 200.100000 56.240000 ;
      RECT 1.000000 54.800000 199.100000 55.780000 ;
      RECT 0.000000 54.600000 200.100000 54.800000 ;
      RECT 197.570000 54.560000 200.100000 54.600000 ;
      RECT 0.000000 54.560000 2.530000 54.600000 ;
      RECT 197.570000 53.580000 199.100000 54.560000 ;
      RECT 1.000000 53.580000 2.530000 54.560000 ;
      RECT 197.570000 53.520000 200.100000 53.580000 ;
      RECT 188.560000 53.520000 195.770000 54.600000 ;
      RECT 143.560000 53.520000 186.760000 54.600000 ;
      RECT 98.560000 53.520000 141.760000 54.600000 ;
      RECT 53.560000 53.520000 96.760000 54.600000 ;
      RECT 8.560000 53.520000 51.760000 54.600000 ;
      RECT 4.330000 53.520000 6.760000 54.600000 ;
      RECT 0.000000 53.520000 2.530000 53.580000 ;
      RECT 0.000000 53.340000 200.100000 53.520000 ;
      RECT 1.000000 52.360000 199.100000 53.340000 ;
      RECT 0.000000 51.880000 200.100000 52.360000 ;
      RECT 199.370000 51.510000 200.100000 51.880000 ;
      RECT 0.000000 51.510000 0.730000 51.880000 ;
      RECT 186.560000 50.800000 197.570000 51.880000 ;
      RECT 141.560000 50.800000 184.760000 51.880000 ;
      RECT 96.560000 50.800000 139.760000 51.880000 ;
      RECT 51.560000 50.800000 94.760000 51.880000 ;
      RECT 6.560000 50.800000 49.760000 51.880000 ;
      RECT 2.530000 50.800000 4.595000 51.880000 ;
      RECT 1.000000 50.530000 199.100000 50.800000 ;
      RECT 0.000000 50.290000 200.100000 50.530000 ;
      RECT 1.000000 49.310000 199.100000 50.290000 ;
      RECT 0.000000 49.160000 200.100000 49.310000 ;
      RECT 197.570000 48.460000 200.100000 49.160000 ;
      RECT 0.000000 48.460000 2.530000 49.160000 ;
      RECT 197.570000 48.080000 199.100000 48.460000 ;
      RECT 188.560000 48.080000 195.770000 49.160000 ;
      RECT 143.560000 48.080000 186.760000 49.160000 ;
      RECT 98.560000 48.080000 141.760000 49.160000 ;
      RECT 53.560000 48.080000 96.760000 49.160000 ;
      RECT 8.560000 48.080000 51.760000 49.160000 ;
      RECT 4.330000 48.080000 6.760000 49.160000 ;
      RECT 1.000000 48.080000 2.530000 48.460000 ;
      RECT 1.000000 47.480000 199.100000 48.080000 ;
      RECT 0.000000 47.240000 200.100000 47.480000 ;
      RECT 1.000000 46.440000 199.100000 47.240000 ;
      RECT 199.370000 45.410000 200.100000 46.260000 ;
      RECT 0.000000 45.410000 0.730000 46.260000 ;
      RECT 186.560000 45.360000 197.570000 46.440000 ;
      RECT 141.560000 45.360000 184.760000 46.440000 ;
      RECT 96.560000 45.360000 139.760000 46.440000 ;
      RECT 51.560000 45.360000 94.760000 46.440000 ;
      RECT 6.560000 45.360000 49.760000 46.440000 ;
      RECT 2.530000 45.360000 4.595000 46.440000 ;
      RECT 1.000000 44.430000 199.100000 45.360000 ;
      RECT 0.000000 44.190000 200.100000 44.430000 ;
      RECT 1.000000 43.720000 199.100000 44.190000 ;
      RECT 197.570000 43.210000 199.100000 43.720000 ;
      RECT 1.000000 43.210000 2.530000 43.720000 ;
      RECT 197.570000 42.970000 200.100000 43.210000 ;
      RECT 0.000000 42.970000 2.530000 43.210000 ;
      RECT 197.570000 42.640000 199.100000 42.970000 ;
      RECT 188.560000 42.640000 195.770000 43.720000 ;
      RECT 143.560000 42.640000 186.760000 43.720000 ;
      RECT 98.560000 42.640000 141.760000 43.720000 ;
      RECT 53.560000 42.640000 96.760000 43.720000 ;
      RECT 8.560000 42.640000 51.760000 43.720000 ;
      RECT 4.330000 42.640000 6.760000 43.720000 ;
      RECT 1.000000 42.640000 2.530000 42.970000 ;
      RECT 1.000000 41.990000 199.100000 42.640000 ;
      RECT 0.000000 41.140000 200.100000 41.990000 ;
      RECT 1.000000 41.000000 199.100000 41.140000 ;
      RECT 199.370000 39.920000 200.100000 40.160000 ;
      RECT 186.560000 39.920000 197.570000 41.000000 ;
      RECT 141.560000 39.920000 184.760000 41.000000 ;
      RECT 96.560000 39.920000 139.760000 41.000000 ;
      RECT 51.560000 39.920000 94.760000 41.000000 ;
      RECT 6.560000 39.920000 49.760000 41.000000 ;
      RECT 2.530000 39.920000 4.595000 41.000000 ;
      RECT 0.000000 39.920000 0.730000 40.160000 ;
      RECT 1.000000 38.940000 199.100000 39.920000 ;
      RECT 0.000000 38.280000 200.100000 38.940000 ;
      RECT 197.570000 38.090000 200.100000 38.280000 ;
      RECT 0.000000 38.090000 2.530000 38.280000 ;
      RECT 197.570000 37.200000 199.100000 38.090000 ;
      RECT 188.560000 37.200000 195.770000 38.280000 ;
      RECT 143.560000 37.200000 186.760000 38.280000 ;
      RECT 98.560000 37.200000 141.760000 38.280000 ;
      RECT 53.560000 37.200000 96.760000 38.280000 ;
      RECT 8.560000 37.200000 51.760000 38.280000 ;
      RECT 4.330000 37.200000 6.760000 38.280000 ;
      RECT 1.000000 37.200000 2.530000 38.090000 ;
      RECT 1.000000 37.110000 199.100000 37.200000 ;
      RECT 0.000000 36.870000 200.100000 37.110000 ;
      RECT 1.000000 35.890000 199.100000 36.870000 ;
      RECT 0.000000 35.560000 200.100000 35.890000 ;
      RECT 199.370000 35.040000 200.100000 35.560000 ;
      RECT 0.000000 35.040000 0.730000 35.560000 ;
      RECT 186.560000 34.480000 197.570000 35.560000 ;
      RECT 141.560000 34.480000 184.760000 35.560000 ;
      RECT 96.560000 34.480000 139.760000 35.560000 ;
      RECT 51.560000 34.480000 94.760000 35.560000 ;
      RECT 6.560000 34.480000 49.760000 35.560000 ;
      RECT 2.530000 34.480000 4.595000 35.560000 ;
      RECT 1.000000 34.060000 199.100000 34.480000 ;
      RECT 0.000000 33.820000 200.100000 34.060000 ;
      RECT 1.000000 32.840000 199.100000 33.820000 ;
      RECT 197.570000 31.990000 200.100000 32.840000 ;
      RECT 0.000000 31.990000 2.530000 32.840000 ;
      RECT 197.570000 31.760000 199.100000 31.990000 ;
      RECT 188.560000 31.760000 195.770000 32.840000 ;
      RECT 143.560000 31.760000 186.760000 32.840000 ;
      RECT 98.560000 31.760000 141.760000 32.840000 ;
      RECT 53.560000 31.760000 96.760000 32.840000 ;
      RECT 8.560000 31.760000 51.760000 32.840000 ;
      RECT 4.330000 31.760000 6.760000 32.840000 ;
      RECT 1.000000 31.760000 2.530000 31.990000 ;
      RECT 1.000000 31.010000 199.100000 31.760000 ;
      RECT 0.000000 30.770000 200.100000 31.010000 ;
      RECT 1.000000 30.120000 199.100000 30.770000 ;
      RECT 199.370000 29.550000 200.100000 29.790000 ;
      RECT 0.000000 29.550000 0.730000 29.790000 ;
      RECT 186.560000 29.040000 197.570000 30.120000 ;
      RECT 141.560000 29.040000 184.760000 30.120000 ;
      RECT 96.560000 29.040000 139.760000 30.120000 ;
      RECT 51.560000 29.040000 94.760000 30.120000 ;
      RECT 6.560000 29.040000 49.760000 30.120000 ;
      RECT 2.530000 29.040000 4.595000 30.120000 ;
      RECT 1.000000 28.570000 199.100000 29.040000 ;
      RECT 0.000000 27.720000 200.100000 28.570000 ;
      RECT 1.000000 27.400000 199.100000 27.720000 ;
      RECT 197.570000 26.740000 199.100000 27.400000 ;
      RECT 1.000000 26.740000 2.530000 27.400000 ;
      RECT 197.570000 26.500000 200.100000 26.740000 ;
      RECT 0.000000 26.500000 2.530000 26.740000 ;
      RECT 197.570000 26.320000 199.100000 26.500000 ;
      RECT 188.560000 26.320000 195.770000 27.400000 ;
      RECT 143.560000 26.320000 186.760000 27.400000 ;
      RECT 98.560000 26.320000 141.760000 27.400000 ;
      RECT 53.560000 26.320000 96.760000 27.400000 ;
      RECT 8.560000 26.320000 51.760000 27.400000 ;
      RECT 4.330000 26.320000 6.760000 27.400000 ;
      RECT 1.000000 26.320000 2.530000 26.500000 ;
      RECT 1.000000 25.520000 199.100000 26.320000 ;
      RECT 0.000000 24.680000 200.100000 25.520000 ;
      RECT 199.370000 24.670000 200.100000 24.680000 ;
      RECT 0.000000 24.670000 0.730000 24.680000 ;
      RECT 199.370000 23.600000 200.100000 23.690000 ;
      RECT 186.560000 23.600000 197.570000 24.680000 ;
      RECT 141.560000 23.600000 184.760000 24.680000 ;
      RECT 96.560000 23.600000 139.760000 24.680000 ;
      RECT 51.560000 23.600000 94.760000 24.680000 ;
      RECT 6.560000 23.600000 49.760000 24.680000 ;
      RECT 2.530000 23.600000 4.595000 24.680000 ;
      RECT 0.000000 23.600000 0.730000 23.690000 ;
      RECT 0.000000 23.450000 200.100000 23.600000 ;
      RECT 1.000000 22.470000 199.100000 23.450000 ;
      RECT 0.000000 21.960000 200.100000 22.470000 ;
      RECT 197.570000 21.620000 200.100000 21.960000 ;
      RECT 0.000000 21.620000 2.530000 21.960000 ;
      RECT 197.570000 20.880000 199.100000 21.620000 ;
      RECT 188.560000 20.880000 195.770000 21.960000 ;
      RECT 143.560000 20.880000 186.760000 21.960000 ;
      RECT 98.560000 20.880000 141.760000 21.960000 ;
      RECT 53.560000 20.880000 96.760000 21.960000 ;
      RECT 8.560000 20.880000 51.760000 21.960000 ;
      RECT 4.330000 20.880000 6.760000 21.960000 ;
      RECT 1.000000 20.880000 2.530000 21.620000 ;
      RECT 1.000000 20.640000 199.100000 20.880000 ;
      RECT 0.000000 20.400000 200.100000 20.640000 ;
      RECT 1.000000 19.420000 199.100000 20.400000 ;
      RECT 0.000000 19.240000 200.100000 19.420000 ;
      RECT 199.370000 18.570000 200.100000 19.240000 ;
      RECT 0.000000 18.570000 0.730000 19.240000 ;
      RECT 186.560000 18.160000 197.570000 19.240000 ;
      RECT 141.560000 18.160000 184.760000 19.240000 ;
      RECT 96.560000 18.160000 139.760000 19.240000 ;
      RECT 51.560000 18.160000 94.760000 19.240000 ;
      RECT 6.560000 18.160000 49.760000 19.240000 ;
      RECT 2.530000 18.160000 4.595000 19.240000 ;
      RECT 1.000000 17.590000 199.100000 18.160000 ;
      RECT 0.000000 17.350000 200.100000 17.590000 ;
      RECT 1.000000 16.520000 199.100000 17.350000 ;
      RECT 197.570000 16.370000 199.100000 16.520000 ;
      RECT 1.000000 16.370000 2.530000 16.520000 ;
      RECT 197.570000 16.130000 200.100000 16.370000 ;
      RECT 0.000000 16.130000 2.530000 16.370000 ;
      RECT 197.570000 15.440000 199.100000 16.130000 ;
      RECT 188.560000 15.440000 195.770000 16.520000 ;
      RECT 143.560000 15.440000 186.760000 16.520000 ;
      RECT 98.560000 15.440000 141.760000 16.520000 ;
      RECT 53.560000 15.440000 96.760000 16.520000 ;
      RECT 8.560000 15.440000 51.760000 16.520000 ;
      RECT 4.330000 15.440000 6.760000 16.520000 ;
      RECT 1.000000 15.440000 2.530000 16.130000 ;
      RECT 1.000000 15.150000 199.100000 15.440000 ;
      RECT 0.000000 14.300000 200.100000 15.150000 ;
      RECT 1.000000 13.800000 199.100000 14.300000 ;
      RECT 199.370000 13.080000 200.100000 13.320000 ;
      RECT 0.000000 13.080000 0.730000 13.320000 ;
      RECT 186.560000 12.720000 197.570000 13.800000 ;
      RECT 141.560000 12.720000 184.760000 13.800000 ;
      RECT 96.560000 12.720000 139.760000 13.800000 ;
      RECT 51.560000 12.720000 94.760000 13.800000 ;
      RECT 6.560000 12.720000 49.760000 13.800000 ;
      RECT 2.530000 12.720000 4.595000 13.800000 ;
      RECT 1.000000 12.100000 199.100000 12.720000 ;
      RECT 0.000000 11.250000 200.100000 12.100000 ;
      RECT 1.000000 11.080000 199.100000 11.250000 ;
      RECT 197.570000 10.270000 199.100000 11.080000 ;
      RECT 1.000000 10.270000 2.530000 11.080000 ;
      RECT 197.570000 10.030000 200.100000 10.270000 ;
      RECT 0.000000 10.030000 2.530000 10.270000 ;
      RECT 197.570000 10.000000 199.100000 10.030000 ;
      RECT 188.560000 10.000000 195.770000 11.080000 ;
      RECT 143.560000 10.000000 186.760000 11.080000 ;
      RECT 98.560000 10.000000 141.760000 11.080000 ;
      RECT 53.560000 10.000000 96.760000 11.080000 ;
      RECT 8.560000 10.000000 51.760000 11.080000 ;
      RECT 4.330000 10.000000 6.760000 11.080000 ;
      RECT 1.000000 10.000000 2.530000 10.030000 ;
      RECT 1.000000 9.050000 199.100000 10.000000 ;
      RECT 0.000000 8.360000 200.100000 9.050000 ;
      RECT 199.370000 8.200000 200.100000 8.360000 ;
      RECT 0.000000 8.200000 0.730000 8.360000 ;
      RECT 186.560000 7.280000 197.570000 8.360000 ;
      RECT 141.560000 7.280000 184.760000 8.360000 ;
      RECT 96.560000 7.280000 139.760000 8.360000 ;
      RECT 51.560000 7.280000 94.760000 8.360000 ;
      RECT 6.560000 7.280000 49.760000 8.360000 ;
      RECT 2.530000 7.280000 4.595000 8.360000 ;
      RECT 1.000000 7.220000 199.100000 7.280000 ;
      RECT 0.000000 6.980000 200.100000 7.220000 ;
      RECT 1.000000 6.000000 199.100000 6.980000 ;
      RECT 0.000000 5.760000 200.100000 6.000000 ;
      RECT 1.000000 5.640000 199.100000 5.760000 ;
      RECT 197.570000 4.780000 199.100000 5.640000 ;
      RECT 1.000000 4.780000 2.530000 5.640000 ;
      RECT 197.570000 4.560000 200.100000 4.780000 ;
      RECT 188.560000 4.560000 195.770000 5.640000 ;
      RECT 143.560000 4.560000 186.760000 5.640000 ;
      RECT 98.560000 4.560000 141.760000 5.640000 ;
      RECT 53.560000 4.560000 96.760000 5.640000 ;
      RECT 8.560000 4.560000 51.760000 5.640000 ;
      RECT 4.330000 4.560000 6.760000 5.640000 ;
      RECT 0.000000 4.560000 2.530000 4.780000 ;
      RECT 0.000000 4.350000 200.100000 4.560000 ;
      RECT 0.000000 0.000000 200.100000 0.750000 ;
    LAYER met4 ;
      RECT 4.330000 198.320000 195.770000 200.260000 ;
      RECT 186.560000 196.520000 195.770000 198.320000 ;
      RECT 141.560000 196.520000 184.760000 198.320000 ;
      RECT 96.560000 196.520000 139.760000 198.320000 ;
      RECT 51.560000 196.520000 94.760000 198.320000 ;
      RECT 6.560000 196.520000 49.760000 198.320000 ;
      RECT 4.330000 193.320000 4.760000 198.320000 ;
      RECT 4.330000 192.240000 4.595000 193.320000 ;
      RECT 4.330000 187.880000 4.760000 192.240000 ;
      RECT 4.330000 186.800000 4.595000 187.880000 ;
      RECT 4.330000 182.440000 4.760000 186.800000 ;
      RECT 4.330000 181.360000 4.595000 182.440000 ;
      RECT 4.330000 177.000000 4.760000 181.360000 ;
      RECT 4.330000 175.920000 4.595000 177.000000 ;
      RECT 4.330000 171.560000 4.760000 175.920000 ;
      RECT 4.330000 170.480000 4.595000 171.560000 ;
      RECT 4.330000 166.120000 4.760000 170.480000 ;
      RECT 4.330000 165.040000 4.595000 166.120000 ;
      RECT 4.330000 160.680000 4.760000 165.040000 ;
      RECT 4.330000 159.600000 4.595000 160.680000 ;
      RECT 4.330000 155.240000 4.760000 159.600000 ;
      RECT 4.330000 154.160000 4.595000 155.240000 ;
      RECT 4.330000 149.800000 4.760000 154.160000 ;
      RECT 4.330000 148.720000 4.595000 149.800000 ;
      RECT 4.330000 144.360000 4.760000 148.720000 ;
      RECT 4.330000 143.280000 4.595000 144.360000 ;
      RECT 4.330000 138.920000 4.760000 143.280000 ;
      RECT 4.330000 137.840000 4.595000 138.920000 ;
      RECT 4.330000 133.480000 4.760000 137.840000 ;
      RECT 4.330000 132.400000 4.595000 133.480000 ;
      RECT 4.330000 128.040000 4.760000 132.400000 ;
      RECT 4.330000 126.960000 4.595000 128.040000 ;
      RECT 4.330000 122.600000 4.760000 126.960000 ;
      RECT 4.330000 121.520000 4.595000 122.600000 ;
      RECT 4.330000 117.160000 4.760000 121.520000 ;
      RECT 4.330000 116.080000 4.595000 117.160000 ;
      RECT 4.330000 111.720000 4.760000 116.080000 ;
      RECT 4.330000 110.640000 4.595000 111.720000 ;
      RECT 4.330000 106.280000 4.760000 110.640000 ;
      RECT 4.330000 105.200000 4.595000 106.280000 ;
      RECT 4.330000 100.840000 4.760000 105.200000 ;
      RECT 4.330000 99.760000 4.595000 100.840000 ;
      RECT 4.330000 95.400000 4.760000 99.760000 ;
      RECT 4.330000 94.320000 4.595000 95.400000 ;
      RECT 4.330000 89.960000 4.760000 94.320000 ;
      RECT 4.330000 88.880000 4.595000 89.960000 ;
      RECT 4.330000 84.520000 4.760000 88.880000 ;
      RECT 4.330000 83.440000 4.595000 84.520000 ;
      RECT 4.330000 79.080000 4.760000 83.440000 ;
      RECT 4.330000 78.000000 4.595000 79.080000 ;
      RECT 4.330000 73.640000 4.760000 78.000000 ;
      RECT 4.330000 72.560000 4.595000 73.640000 ;
      RECT 4.330000 68.200000 4.760000 72.560000 ;
      RECT 4.330000 67.120000 4.595000 68.200000 ;
      RECT 4.330000 62.760000 4.760000 67.120000 ;
      RECT 4.330000 61.680000 4.595000 62.760000 ;
      RECT 4.330000 57.320000 4.760000 61.680000 ;
      RECT 4.330000 56.240000 4.595000 57.320000 ;
      RECT 4.330000 51.880000 4.760000 56.240000 ;
      RECT 4.330000 50.800000 4.595000 51.880000 ;
      RECT 4.330000 46.440000 4.760000 50.800000 ;
      RECT 4.330000 45.360000 4.595000 46.440000 ;
      RECT 4.330000 41.000000 4.760000 45.360000 ;
      RECT 4.330000 39.920000 4.595000 41.000000 ;
      RECT 4.330000 35.560000 4.760000 39.920000 ;
      RECT 4.330000 34.480000 4.595000 35.560000 ;
      RECT 4.330000 30.120000 4.760000 34.480000 ;
      RECT 4.330000 29.040000 4.595000 30.120000 ;
      RECT 4.330000 24.680000 4.760000 29.040000 ;
      RECT 4.330000 23.600000 4.595000 24.680000 ;
      RECT 4.330000 19.240000 4.760000 23.600000 ;
      RECT 4.330000 18.160000 4.595000 19.240000 ;
      RECT 4.330000 13.800000 4.760000 18.160000 ;
      RECT 4.330000 12.720000 4.595000 13.800000 ;
      RECT 4.330000 8.360000 4.760000 12.720000 ;
      RECT 4.330000 7.280000 4.595000 8.360000 ;
      RECT 188.560000 2.550000 195.770000 196.520000 ;
      RECT 186.560000 2.550000 186.760000 196.520000 ;
      RECT 143.560000 2.550000 184.760000 196.520000 ;
      RECT 141.560000 2.550000 141.760000 196.520000 ;
      RECT 98.560000 2.550000 139.760000 196.520000 ;
      RECT 96.560000 2.550000 96.760000 196.520000 ;
      RECT 53.560000 2.550000 94.760000 196.520000 ;
      RECT 51.560000 2.550000 51.760000 196.520000 ;
      RECT 8.560000 2.550000 49.760000 196.520000 ;
      RECT 6.560000 2.550000 6.760000 196.520000 ;
      RECT 186.560000 0.750000 195.770000 2.550000 ;
      RECT 141.560000 0.750000 184.760000 2.550000 ;
      RECT 96.560000 0.750000 139.760000 2.550000 ;
      RECT 51.560000 0.750000 94.760000 2.550000 ;
      RECT 6.560000 0.750000 49.760000 2.550000 ;
      RECT 4.330000 0.750000 4.760000 7.280000 ;
      RECT 199.370000 0.000000 200.100000 200.260000 ;
      RECT 4.330000 0.000000 195.770000 0.750000 ;
      RECT 0.000000 0.000000 0.730000 200.260000 ;
  END
END LUT4AB

END LIBRARY
