##
## LEF for PtnCells ;
## created by Innovus v19.11-s128_1 on Tue Nov 23 23:01:49 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO N_term_single
  CLASS BLOCK ;
  SIZE 200.100000 BY 30.260000 ;
  FOREIGN N_term_single 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.912 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.452 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.68323 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 27.035 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 9.240000 0.000000 9.620000 0.700000 ;
    END
  END N1END[3]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.955 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.94997 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.0774 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 7.860000 0.000000 8.240000 0.700000 ;
    END
  END N1END[2]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.129 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.537 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.56357 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.4431 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 6.480000 0.000000 6.860000 0.700000 ;
    END
  END N1END[1]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4482 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.133 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.63697 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.8101 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 0.000000 5.480000 0.700000 ;
    END
  END N1END[0]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0602 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.075 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.02505 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.58519 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 21.660000 0.000000 22.040000 0.700000 ;
    END
  END N2MID[7]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.129 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.537 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.20741 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.6559 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 19.820000 0.000000 20.200000 0.700000 ;
    END
  END N2MID[6]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2299 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.5008 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 8.03879 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 42.0229 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 18.440000 0.000000 18.820000 0.700000 ;
    END
  END N2MID[5]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.0048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.496 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 9.10545 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 47.4815 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 17.060000 0.000000 17.440000 0.700000 ;
    END
  END N2MID[4]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8029 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.5588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.784 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 18.04 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 94.1077 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 15.680000 0.000000 16.060000 0.700000 ;
    END
  END N2MID[3]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6526 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.155 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.7429 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.3333 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 13.840000 0.000000 14.220000 0.700000 ;
    END
  END N2MID[2]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6569 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.7328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 19.2812 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 101.832 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 12.460000 0.000000 12.840000 0.700000 ;
    END
  END N2MID[1]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.846 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.26613 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.936 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 11.080000 0.000000 11.460000 0.700000 ;
    END
  END N2MID[0]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7478 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.631 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.38034 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.5205 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 33.620000 0.000000 34.000000 0.700000 ;
    END
  END N2END[7]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.441 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.47805 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.2101 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 32.240000 0.000000 32.620000 0.700000 ;
    END
  END N2END[6]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4861 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.1908 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.488 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 11.4671 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 59.2822 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 30.860000 0.000000 31.240000 0.700000 ;
    END
  END N2END[5]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7482 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.633 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.02963 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.767 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 29.020000 0.000000 29.400000 0.700000 ;
    END
  END N2END[4]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.367 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.727 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.18155 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.5266 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 27.640000 0.000000 28.020000 0.700000 ;
    END
  END N2END[3]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.0528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.752 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 10.5232 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 54.501 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 26.260000 0.000000 26.640000 0.700000 ;
    END
  END N2END[2]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8698 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.123 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.76721 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.602 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 24.420000 0.000000 24.800000 0.700000 ;
    END
  END N2END[1]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2242 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.013 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.61104 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 16.6741 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 23.040000 0.000000 23.420000 0.700000 ;
    END
  END N2END[0]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4861 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.2848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.656 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 20.8069 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 109.615 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 58.000000 0.000000 58.380000 0.700000 ;
    END
  END N4END[15]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0602 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.075 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.84646 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.6923 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 56.620000 0.000000 57.000000 0.700000 ;
    END
  END N4END[14]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7482 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.633 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.18687 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 28.262 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 54.780000 0.000000 55.160000 0.700000 ;
    END
  END N4END[13]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5222 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.385 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.02936 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.6067 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 53.400000 0.000000 53.780000 0.700000 ;
    END
  END N4END[12]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.2258 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.008 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 20.2423 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 106.316 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 52.020000 0.000000 52.400000 0.700000 ;
    END
  END N4END[11]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.703 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.407 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.07508 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.2983 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 50.180000 0.000000 50.560000 0.700000 ;
    END
  END N4END[10]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.967 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.14316 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.1758 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 48.800000 0.000000 49.180000 0.700000 ;
    END
  END N4END[9]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.829 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.037 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.15583 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.398 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 47.420000 0.000000 47.800000 0.700000 ;
    END
  END N4END[8]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9493 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.6748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.736 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 12.9572 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 67.8478 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 45.580000 0.000000 45.960000 0.700000 ;
    END
  END N4END[7]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.129 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.537 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.60882 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.6694 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 44.200000 0.000000 44.580000 0.700000 ;
    END
  END N4END[6]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.837 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.82397 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.67071 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 42.820000 0.000000 43.200000 0.700000 ;
    END
  END N4END[5]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.115 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.467 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.34505 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.3441 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 41.440000 0.000000 41.820000 0.700000 ;
    END
  END N4END[4]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0381 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.4428 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.832 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 17.9244 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 94.3758 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 39.600000 0.000000 39.980000 0.700000 ;
    END
  END N4END[3]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.6538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.624 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 21.4453 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 112.972 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 38.220000 0.000000 38.600000 0.700000 ;
    END
  END N4END[2]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7054 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.183 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.82424 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 12.4222 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 36.840000 0.000000 37.220000 0.700000 ;
    END
  END N4END[1]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.837 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.06465 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.78316 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 35.000000 0.000000 35.380000 0.700000 ;
    END
  END N4END[0]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.502 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.0031 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.56633 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 82.380000 0.000000 82.760000 0.700000 ;
    END
  END NN4END[15]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.441 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.02249 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.7313 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 80.540000 0.000000 80.920000 0.700000 ;
    END
  END NN4END[14]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3458 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.503 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.27273 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 9.91448 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 79.160000 0.000000 79.540000 0.700000 ;
    END
  END NN4END[13]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.441 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.979 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.23508 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.3441 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 77.780000 0.000000 78.160000 0.700000 ;
    END
  END NN4END[12]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0336 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.942 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.85226 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.81212 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 75.940000 0.000000 76.320000 0.700000 ;
    END
  END NN4END[11]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.367 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.727 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.74788 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.3582 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 74.560000 0.000000 74.940000 0.700000 ;
    END
  END NN4END[10]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6102 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.707 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.62882 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 11.536 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 73.180000 0.000000 73.560000 0.700000 ;
    END
  END NN4END[9]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4479 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.0785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.3568 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.04 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 30.4648 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 160.63 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 71.800000 0.000000 72.180000 0.700000 ;
    END
  END NN4END[8]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5358 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.453 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.94263 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.1731 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 69.960000 0.000000 70.340000 0.700000 ;
    END
  END NN4END[7]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.569 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.619 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.26694 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.8855 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 68.580000 0.000000 68.960000 0.700000 ;
    END
  END NN4END[6]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6569 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.1928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 118.832 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 30.6341 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 162.392 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 67.200000 0.000000 67.580000 0.700000 ;
    END
  END NN4END[5]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9382 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.583 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 15.5143 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 76.1906 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 65.360000 0.000000 65.740000 0.700000 ;
    END
  END NN4END[4]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.441 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 10.1074 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 48.0572 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 63.980000 0.000000 64.360000 0.700000 ;
    END
  END NN4END[3]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1445 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.6308 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.168 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 23.7779 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 125.523 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 62.600000 0.000000 62.980000 0.700000 ;
    END
  END NN4END[2]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.997 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.759 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.19017 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.5017 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 60.760000 0.000000 61.140000 0.700000 ;
    END
  END NN4END[1]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.92054 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.20808 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 59.380000 0.000000 59.760000 0.700000 ;
    END
  END NN4END[0]
  PIN Ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.260000 0.000000 164.640000 0.700000 ;
    END
  END Ci
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6208 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.943 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.1488 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.264 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 88.360000 0.000000 88.740000 0.700000 ;
    END
  END S1BEG[3]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.2042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.795 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 86.520000 0.000000 86.900000 0.700000 ;
    END
  END S1BEG[2]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0142 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.845 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 85.140000 0.000000 85.520000 0.700000 ;
    END
  END S1BEG[1]
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2316 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.997 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.2058 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.568 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 83.760000 0.000000 84.140000 0.700000 ;
    END
  END S1BEG[0]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.4648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.616 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 112.740000 0.000000 113.120000 0.700000 ;
    END
  END S2BEG[7]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.0508 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.408 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 110.900000 0.000000 111.280000 0.700000 ;
    END
  END S2BEG[6]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.6354 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.951 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 109.520000 0.000000 109.900000 0.700000 ;
    END
  END S2BEG[5]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8029 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.3058 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.768 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 108.140000 0.000000 108.520000 0.700000 ;
    END
  END S2BEG[4]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7671 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.1288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 107.824 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 106.300000 0.000000 106.680000 0.700000 ;
    END
  END S2BEG[3]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2795 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.2365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.7118 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.6 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 104.920000 0.000000 105.300000 0.700000 ;
    END
  END S2BEG[2]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8378 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.963 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 103.540000 0.000000 103.920000 0.700000 ;
    END
  END S2BEG[1]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.5708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.848 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 101.700000 0.000000 102.080000 0.700000 ;
    END
  END S2BEG[0]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.5062 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.305 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 100.320000 0.000000 100.700000 0.700000 ;
    END
  END S2BEGb[7]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.059 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 98.940000 0.000000 99.320000 0.700000 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9246 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.515 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 97.560000 0.000000 97.940000 0.700000 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.441 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.979 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 95.720000 0.000000 96.100000 0.700000 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.0166 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.857 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 94.340000 0.000000 94.720000 0.700000 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0591 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.1345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.3608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 92.960000 0.000000 93.340000 0.700000 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.7898 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.016 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 91.120000 0.000000 91.500000 0.700000 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.2046 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.797 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 89.740000 0.000000 90.120000 0.700000 ;
    END
  END S2BEGb[0]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.431 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 136.660000 0.000000 137.040000 0.700000 ;
    END
  END S4BEG[15]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.837 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 135.280000 0.000000 135.660000 0.700000 ;
    END
  END S4BEG[14]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1025 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.8828 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.512 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 133.900000 0.000000 134.280000 0.700000 ;
    END
  END S4BEG[13]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5963 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.9416 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.296 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 132.060000 0.000000 132.440000 0.700000 ;
    END
  END S4BEG[12]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0595 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.0185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.2608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.528 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 130.680000 0.000000 131.060000 0.700000 ;
    END
  END S4BEG[11]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.837 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 129.300000 0.000000 129.680000 0.700000 ;
    END
  END S4BEG[10]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1979 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.8285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.6468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 115.92 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 127.460000 0.000000 127.840000 0.700000 ;
    END
  END S4BEG[9]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.8458 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.648 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 126.080000 0.000000 126.460000 0.700000 ;
    END
  END S4BEG[8]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.4136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.842 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 124.700000 0.000000 125.080000 0.700000 ;
    END
  END S4BEG[7]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8277 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.9775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.1228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.792 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 123.320000 0.000000 123.700000 0.700000 ;
    END
  END S4BEG[6]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3314 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.431 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 121.480000 0.000000 121.860000 0.700000 ;
    END
  END S4BEG[5]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.5458 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.048 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 120.100000 0.000000 120.480000 0.700000 ;
    END
  END S4BEG[4]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.741 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 118.720000 0.000000 119.100000 0.700000 ;
    END
  END S4BEG[3]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.837 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 116.880000 0.000000 117.260000 0.700000 ;
    END
  END S4BEG[2]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.823 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 115.500000 0.000000 115.880000 0.700000 ;
    END
  END S4BEG[1]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6526 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.155 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 114.120000 0.000000 114.500000 0.700000 ;
    END
  END S4BEG[0]
  PIN SS4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.502 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 161.040000 0.000000 161.420000 0.700000 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5574 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.679 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 159.660000 0.000000 160.040000 0.700000 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.599 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.820000 0.000000 158.200000 0.700000 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5715 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.6828 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.112 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 156.440000 0.000000 156.820000 0.700000 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9382 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.583 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 155.060000 0.000000 155.440000 0.700000 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7646 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.715 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 153.680000 0.000000 154.060000 0.700000 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.88 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 151.840000 0.000000 152.220000 0.700000 ;
    END
  END SS4BEG[9]
  PIN SS4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.784 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.460000 0.000000 150.840000 0.700000 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8434 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.109 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 149.080000 0.000000 149.460000 0.700000 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7768 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.28 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 147.240000 0.000000 147.620000 0.700000 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9174 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.361 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 145.860000 0.000000 146.240000 0.700000 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.077 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.159 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 144.480000 0.000000 144.860000 0.700000 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4006 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.895 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 142.640000 0.000000 143.020000 0.700000 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3626 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.587 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 141.260000 0.000000 141.640000 0.700000 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.717 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.477 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 139.880000 0.000000 140.260000 0.700000 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.871 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 138.500000 0.000000 138.880000 0.700000 ;
    END
  END SS4BEG[0]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2299 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.5368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.152 LAYER met3  ;
    ANTENNAMAXAREACAR 8.05831 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 41.3385 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.0793403 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 162.420000 0.000000 162.800000 0.700000 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3218 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.501 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 29.560000 5.480000 30.260000 ;
    END
  END UserCLKo
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7474 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.629 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.83475 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.7926 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 194.160000 0.000000 194.540000 0.700000 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2714 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.249 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.92424 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 16.9488 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 192.780000 0.000000 193.160000 0.700000 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6522 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.153 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.72034 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.8242 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 191.400000 0.000000 191.780000 0.700000 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8426 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.105 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.65805 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.9091 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 190.020000 0.000000 190.400000 0.700000 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.308 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.04909 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.7118 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 188.180000 0.000000 188.560000 0.700000 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9978 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.763 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.49764 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.0391 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 186.800000 0.000000 187.180000 0.700000 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.035 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.73333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 47.2855 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 185.420000 0.000000 185.800000 0.700000 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8858 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.203 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.3468 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.2848 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 183.580000 0.000000 183.960000 0.700000 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.9388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.144 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 18.5624 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 97.4303 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 182.200000 0.000000 182.580000 0.700000 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8214 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.881 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.26007 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.8512 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 180.820000 0.000000 181.200000 0.700000 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7396 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.58 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.83293 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 36.3737 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 179.440000 0.000000 179.820000 0.700000 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8214 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.881 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.26007 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.8512 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 177.600000 0.000000 177.980000 0.700000 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7671 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.4328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.112 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 17.6828 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 90.1293 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 176.220000 0.000000 176.600000 0.700000 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8029 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.5768 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.88 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 29.6544 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 156.319 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 174.840000 0.000000 175.220000 0.700000 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1483 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.5805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.0228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 22.101 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 116.434 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 173.000000 0.000000 173.380000 0.700000 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4255 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.9665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.1968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.52 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 26.1017 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 137.686 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 171.620000 0.000000 172.000000 0.700000 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0114 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.831 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.19017 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.4108 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 170.240000 0.000000 170.620000 0.700000 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4878 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.213 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.31152 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.0175 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 168.400000 0.000000 168.780000 0.700000 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.997 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.759 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.86451 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.7825 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 167.020000 0.000000 167.400000 0.700000 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1731 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.7045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.5448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.376 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 36.5485 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 191.638 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 165.640000 0.000000 166.020000 0.700000 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3194 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.489 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 194.620000 29.560000 195.000000 30.260000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.359 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 184.960000 29.560000 185.340000 30.260000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.217 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 175.300000 29.560000 175.680000 30.260000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4006 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.895 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 166.100000 29.560000 166.480000 30.260000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.251 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 156.440000 29.560000 156.820000 30.260000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4622 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.203 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 147.240000 29.560000 147.620000 30.260000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.251 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 137.580000 29.560000 137.960000 30.260000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.392 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 127.920000 29.560000 128.300000 30.260000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.665 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.099 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 118.720000 29.560000 119.100000 30.260000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5362 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.455 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 109.060000 29.560000 109.440000 30.260000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.591 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.847 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.400000 29.560000 99.780000 30.260000 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.272 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 90.200000 29.560000 90.580000 30.260000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.217 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 80.540000 29.560000 80.920000 30.260000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.441 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.979 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 71.340000 29.560000 71.720000 30.260000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.154 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 61.680000 29.560000 62.060000 30.260000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7455 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.5248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.936 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 52.480000 29.560000 52.860000 30.260000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1764 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.656 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 42.820000 29.560000 43.200000 30.260000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.217 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 33.160000 29.560000 33.540000 30.260000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.916 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 23.960000 29.560000 24.340000 30.260000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.217 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 14.300000 29.560000 14.680000 30.260000 ;
    END
  END FrameStrobe_O[0]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 198.900000 25.700000 200.100000 26.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 25.700000 1.200000 26.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.900000 2.850000 200.100000 4.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 1.200000 4.050000 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.070000 29.060000 197.270000 30.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.070000 0.000000 197.270000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 29.060000 4.030000 30.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 0.000000 4.030000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 200.100000 4.050000 ;
        RECT 0.000000 25.700000 200.100000 26.900000 ;
        RECT 7.060000 4.860000 8.260000 5.340000 ;
        RECT 2.830000 4.860000 4.030000 5.340000 ;
        RECT 7.060000 10.300000 8.260000 10.780000 ;
        RECT 2.830000 10.300000 4.030000 10.780000 ;
        RECT 52.060000 10.300000 53.260000 10.780000 ;
        RECT 97.060000 10.300000 98.260000 10.780000 ;
        RECT 97.060000 4.860000 98.260000 5.340000 ;
        RECT 52.060000 4.860000 53.260000 5.340000 ;
        RECT 142.060000 10.300000 143.260000 10.780000 ;
        RECT 142.060000 4.860000 143.260000 5.340000 ;
        RECT 187.060000 4.860000 188.260000 5.340000 ;
        RECT 187.060000 10.300000 188.260000 10.780000 ;
        RECT 196.070000 10.300000 197.270000 10.780000 ;
        RECT 196.070000 4.860000 197.270000 5.340000 ;
        RECT 2.830000 21.180000 4.030000 21.660000 ;
        RECT 7.060000 21.180000 8.260000 21.660000 ;
        RECT 7.060000 15.740000 8.260000 16.220000 ;
        RECT 2.830000 15.740000 4.030000 16.220000 ;
        RECT 52.060000 21.180000 53.260000 21.660000 ;
        RECT 97.060000 21.180000 98.260000 21.660000 ;
        RECT 97.060000 15.740000 98.260000 16.220000 ;
        RECT 52.060000 15.740000 53.260000 16.220000 ;
        RECT 142.060000 21.180000 143.260000 21.660000 ;
        RECT 142.060000 15.740000 143.260000 16.220000 ;
        RECT 187.060000 15.740000 188.260000 16.220000 ;
        RECT 187.060000 21.180000 188.260000 21.660000 ;
        RECT 196.070000 21.180000 197.270000 21.660000 ;
        RECT 196.070000 15.740000 197.270000 16.220000 ;
      LAYER met4 ;
        RECT 187.060000 2.850000 188.260000 26.900000 ;
        RECT 142.060000 2.850000 143.260000 26.900000 ;
        RECT 97.060000 2.850000 98.260000 26.900000 ;
        RECT 52.060000 2.850000 53.260000 26.900000 ;
        RECT 7.060000 2.850000 8.260000 26.900000 ;
        RECT 196.070000 0.000000 197.270000 30.260000 ;
        RECT 2.830000 0.000000 4.030000 30.260000 ;
    END
# end of P/G power stripe data as pin

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 198.900000 27.500000 200.100000 28.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 27.500000 1.200000 28.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.900000 1.050000 200.100000 2.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 1.200000 2.250000 ;
    END
    PORT
      LAYER met4 ;
        RECT 197.870000 29.060000 199.070000 30.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 197.870000 0.000000 199.070000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 29.060000 2.230000 30.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 0.000000 2.230000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 200.100000 2.250000 ;
        RECT 0.000000 27.500000 200.100000 28.700000 ;
        RECT 1.030000 7.580000 2.230000 8.060000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 1.030000 13.020000 2.230000 13.500000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 50.060000 13.020000 51.260000 13.500000 ;
        RECT 95.060000 13.020000 96.260000 13.500000 ;
        RECT 50.060000 7.580000 51.260000 8.060000 ;
        RECT 95.060000 7.580000 96.260000 8.060000 ;
        RECT 140.060000 13.020000 141.260000 13.500000 ;
        RECT 140.060000 7.580000 141.260000 8.060000 ;
        RECT 185.060000 7.580000 186.260000 8.060000 ;
        RECT 185.060000 13.020000 186.260000 13.500000 ;
        RECT 197.870000 7.580000 199.070000 8.060000 ;
        RECT 197.870000 13.020000 199.070000 13.500000 ;
        RECT 1.030000 18.460000 2.230000 18.940000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 1.030000 23.900000 2.230000 24.380000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
        RECT 50.060000 23.900000 51.260000 24.380000 ;
        RECT 95.060000 23.900000 96.260000 24.380000 ;
        RECT 50.060000 18.460000 51.260000 18.940000 ;
        RECT 95.060000 18.460000 96.260000 18.940000 ;
        RECT 140.060000 23.900000 141.260000 24.380000 ;
        RECT 140.060000 18.460000 141.260000 18.940000 ;
        RECT 185.060000 18.460000 186.260000 18.940000 ;
        RECT 185.060000 23.900000 186.260000 24.380000 ;
        RECT 197.870000 18.460000 199.070000 18.940000 ;
        RECT 197.870000 23.900000 199.070000 24.380000 ;
      LAYER met4 ;
        RECT 185.060000 1.050000 186.260000 28.700000 ;
        RECT 140.060000 1.050000 141.260000 28.700000 ;
        RECT 95.060000 1.050000 96.260000 28.700000 ;
        RECT 50.060000 1.050000 51.260000 28.700000 ;
        RECT 5.060000 1.050000 6.260000 28.700000 ;
        RECT 197.870000 0.000000 199.070000 30.260000 ;
        RECT 1.030000 0.000000 2.230000 30.260000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
    END
# end of P/G power stripe data as pin

  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 200.100000 30.260000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 200.100000 30.260000 ;
    LAYER met2 ;
      RECT 195.140000 29.420000 200.100000 30.260000 ;
      RECT 185.480000 29.420000 194.480000 30.260000 ;
      RECT 175.820000 29.420000 184.820000 30.260000 ;
      RECT 166.620000 29.420000 175.160000 30.260000 ;
      RECT 156.960000 29.420000 165.960000 30.260000 ;
      RECT 147.760000 29.420000 156.300000 30.260000 ;
      RECT 138.100000 29.420000 147.100000 30.260000 ;
      RECT 128.440000 29.420000 137.440000 30.260000 ;
      RECT 119.240000 29.420000 127.780000 30.260000 ;
      RECT 109.580000 29.420000 118.580000 30.260000 ;
      RECT 99.920000 29.420000 108.920000 30.260000 ;
      RECT 90.720000 29.420000 99.260000 30.260000 ;
      RECT 81.060000 29.420000 90.060000 30.260000 ;
      RECT 71.860000 29.420000 80.400000 30.260000 ;
      RECT 62.200000 29.420000 71.200000 30.260000 ;
      RECT 53.000000 29.420000 61.540000 30.260000 ;
      RECT 43.340000 29.420000 52.340000 30.260000 ;
      RECT 33.680000 29.420000 42.680000 30.260000 ;
      RECT 24.480000 29.420000 33.020000 30.260000 ;
      RECT 14.820000 29.420000 23.820000 30.260000 ;
      RECT 5.620000 29.420000 14.160000 30.260000 ;
      RECT 0.000000 29.420000 4.960000 30.260000 ;
      RECT 0.000000 0.840000 200.100000 29.420000 ;
      RECT 194.680000 0.000000 200.100000 0.840000 ;
      RECT 193.300000 0.000000 194.020000 0.840000 ;
      RECT 191.920000 0.000000 192.640000 0.840000 ;
      RECT 190.540000 0.000000 191.260000 0.840000 ;
      RECT 188.700000 0.000000 189.880000 0.840000 ;
      RECT 187.320000 0.000000 188.040000 0.840000 ;
      RECT 185.940000 0.000000 186.660000 0.840000 ;
      RECT 184.100000 0.000000 185.280000 0.840000 ;
      RECT 182.720000 0.000000 183.440000 0.840000 ;
      RECT 181.340000 0.000000 182.060000 0.840000 ;
      RECT 179.960000 0.000000 180.680000 0.840000 ;
      RECT 178.120000 0.000000 179.300000 0.840000 ;
      RECT 176.740000 0.000000 177.460000 0.840000 ;
      RECT 175.360000 0.000000 176.080000 0.840000 ;
      RECT 173.520000 0.000000 174.700000 0.840000 ;
      RECT 172.140000 0.000000 172.860000 0.840000 ;
      RECT 170.760000 0.000000 171.480000 0.840000 ;
      RECT 168.920000 0.000000 170.100000 0.840000 ;
      RECT 167.540000 0.000000 168.260000 0.840000 ;
      RECT 166.160000 0.000000 166.880000 0.840000 ;
      RECT 164.780000 0.000000 165.500000 0.840000 ;
      RECT 162.940000 0.000000 164.120000 0.840000 ;
      RECT 161.560000 0.000000 162.280000 0.840000 ;
      RECT 160.180000 0.000000 160.900000 0.840000 ;
      RECT 158.340000 0.000000 159.520000 0.840000 ;
      RECT 156.960000 0.000000 157.680000 0.840000 ;
      RECT 155.580000 0.000000 156.300000 0.840000 ;
      RECT 154.200000 0.000000 154.920000 0.840000 ;
      RECT 152.360000 0.000000 153.540000 0.840000 ;
      RECT 150.980000 0.000000 151.700000 0.840000 ;
      RECT 149.600000 0.000000 150.320000 0.840000 ;
      RECT 147.760000 0.000000 148.940000 0.840000 ;
      RECT 146.380000 0.000000 147.100000 0.840000 ;
      RECT 145.000000 0.000000 145.720000 0.840000 ;
      RECT 143.160000 0.000000 144.340000 0.840000 ;
      RECT 141.780000 0.000000 142.500000 0.840000 ;
      RECT 140.400000 0.000000 141.120000 0.840000 ;
      RECT 139.020000 0.000000 139.740000 0.840000 ;
      RECT 137.180000 0.000000 138.360000 0.840000 ;
      RECT 135.800000 0.000000 136.520000 0.840000 ;
      RECT 134.420000 0.000000 135.140000 0.840000 ;
      RECT 132.580000 0.000000 133.760000 0.840000 ;
      RECT 131.200000 0.000000 131.920000 0.840000 ;
      RECT 129.820000 0.000000 130.540000 0.840000 ;
      RECT 127.980000 0.000000 129.160000 0.840000 ;
      RECT 126.600000 0.000000 127.320000 0.840000 ;
      RECT 125.220000 0.000000 125.940000 0.840000 ;
      RECT 123.840000 0.000000 124.560000 0.840000 ;
      RECT 122.000000 0.000000 123.180000 0.840000 ;
      RECT 120.620000 0.000000 121.340000 0.840000 ;
      RECT 119.240000 0.000000 119.960000 0.840000 ;
      RECT 117.400000 0.000000 118.580000 0.840000 ;
      RECT 116.020000 0.000000 116.740000 0.840000 ;
      RECT 114.640000 0.000000 115.360000 0.840000 ;
      RECT 113.260000 0.000000 113.980000 0.840000 ;
      RECT 111.420000 0.000000 112.600000 0.840000 ;
      RECT 110.040000 0.000000 110.760000 0.840000 ;
      RECT 108.660000 0.000000 109.380000 0.840000 ;
      RECT 106.820000 0.000000 108.000000 0.840000 ;
      RECT 105.440000 0.000000 106.160000 0.840000 ;
      RECT 104.060000 0.000000 104.780000 0.840000 ;
      RECT 102.220000 0.000000 103.400000 0.840000 ;
      RECT 100.840000 0.000000 101.560000 0.840000 ;
      RECT 99.460000 0.000000 100.180000 0.840000 ;
      RECT 98.080000 0.000000 98.800000 0.840000 ;
      RECT 96.240000 0.000000 97.420000 0.840000 ;
      RECT 94.860000 0.000000 95.580000 0.840000 ;
      RECT 93.480000 0.000000 94.200000 0.840000 ;
      RECT 91.640000 0.000000 92.820000 0.840000 ;
      RECT 90.260000 0.000000 90.980000 0.840000 ;
      RECT 88.880000 0.000000 89.600000 0.840000 ;
      RECT 87.040000 0.000000 88.220000 0.840000 ;
      RECT 85.660000 0.000000 86.380000 0.840000 ;
      RECT 84.280000 0.000000 85.000000 0.840000 ;
      RECT 82.900000 0.000000 83.620000 0.840000 ;
      RECT 81.060000 0.000000 82.240000 0.840000 ;
      RECT 79.680000 0.000000 80.400000 0.840000 ;
      RECT 78.300000 0.000000 79.020000 0.840000 ;
      RECT 76.460000 0.000000 77.640000 0.840000 ;
      RECT 75.080000 0.000000 75.800000 0.840000 ;
      RECT 73.700000 0.000000 74.420000 0.840000 ;
      RECT 72.320000 0.000000 73.040000 0.840000 ;
      RECT 70.480000 0.000000 71.660000 0.840000 ;
      RECT 69.100000 0.000000 69.820000 0.840000 ;
      RECT 67.720000 0.000000 68.440000 0.840000 ;
      RECT 65.880000 0.000000 67.060000 0.840000 ;
      RECT 64.500000 0.000000 65.220000 0.840000 ;
      RECT 63.120000 0.000000 63.840000 0.840000 ;
      RECT 61.280000 0.000000 62.460000 0.840000 ;
      RECT 59.900000 0.000000 60.620000 0.840000 ;
      RECT 58.520000 0.000000 59.240000 0.840000 ;
      RECT 57.140000 0.000000 57.860000 0.840000 ;
      RECT 55.300000 0.000000 56.480000 0.840000 ;
      RECT 53.920000 0.000000 54.640000 0.840000 ;
      RECT 52.540000 0.000000 53.260000 0.840000 ;
      RECT 50.700000 0.000000 51.880000 0.840000 ;
      RECT 49.320000 0.000000 50.040000 0.840000 ;
      RECT 47.940000 0.000000 48.660000 0.840000 ;
      RECT 46.100000 0.000000 47.280000 0.840000 ;
      RECT 44.720000 0.000000 45.440000 0.840000 ;
      RECT 43.340000 0.000000 44.060000 0.840000 ;
      RECT 41.960000 0.000000 42.680000 0.840000 ;
      RECT 40.120000 0.000000 41.300000 0.840000 ;
      RECT 38.740000 0.000000 39.460000 0.840000 ;
      RECT 37.360000 0.000000 38.080000 0.840000 ;
      RECT 35.520000 0.000000 36.700000 0.840000 ;
      RECT 34.140000 0.000000 34.860000 0.840000 ;
      RECT 32.760000 0.000000 33.480000 0.840000 ;
      RECT 31.380000 0.000000 32.100000 0.840000 ;
      RECT 29.540000 0.000000 30.720000 0.840000 ;
      RECT 28.160000 0.000000 28.880000 0.840000 ;
      RECT 26.780000 0.000000 27.500000 0.840000 ;
      RECT 24.940000 0.000000 26.120000 0.840000 ;
      RECT 23.560000 0.000000 24.280000 0.840000 ;
      RECT 22.180000 0.000000 22.900000 0.840000 ;
      RECT 20.340000 0.000000 21.520000 0.840000 ;
      RECT 18.960000 0.000000 19.680000 0.840000 ;
      RECT 17.580000 0.000000 18.300000 0.840000 ;
      RECT 16.200000 0.000000 16.920000 0.840000 ;
      RECT 14.360000 0.000000 15.540000 0.840000 ;
      RECT 12.980000 0.000000 13.700000 0.840000 ;
      RECT 11.600000 0.000000 12.320000 0.840000 ;
      RECT 9.760000 0.000000 10.940000 0.840000 ;
      RECT 8.380000 0.000000 9.100000 0.840000 ;
      RECT 7.000000 0.000000 7.720000 0.840000 ;
      RECT 5.620000 0.000000 6.340000 0.840000 ;
      RECT 0.000000 0.000000 4.960000 0.840000 ;
    LAYER met3 ;
      RECT 0.000000 29.000000 200.100000 30.260000 ;
      RECT 0.000000 24.680000 200.100000 25.400000 ;
      RECT 199.370000 23.600000 200.100000 24.680000 ;
      RECT 186.560000 23.600000 197.570000 24.680000 ;
      RECT 141.560000 23.600000 184.760000 24.680000 ;
      RECT 96.560000 23.600000 139.760000 24.680000 ;
      RECT 51.560000 23.600000 94.760000 24.680000 ;
      RECT 6.560000 23.600000 49.760000 24.680000 ;
      RECT 2.530000 23.600000 4.595000 24.680000 ;
      RECT 0.000000 23.600000 0.730000 24.680000 ;
      RECT 0.000000 21.960000 200.100000 23.600000 ;
      RECT 197.570000 20.880000 200.100000 21.960000 ;
      RECT 188.560000 20.880000 195.770000 21.960000 ;
      RECT 143.560000 20.880000 186.760000 21.960000 ;
      RECT 98.560000 20.880000 141.760000 21.960000 ;
      RECT 53.560000 20.880000 96.760000 21.960000 ;
      RECT 8.560000 20.880000 51.760000 21.960000 ;
      RECT 4.330000 20.880000 6.760000 21.960000 ;
      RECT 0.000000 20.880000 2.530000 21.960000 ;
      RECT 0.000000 19.240000 200.100000 20.880000 ;
      RECT 199.370000 18.160000 200.100000 19.240000 ;
      RECT 186.560000 18.160000 197.570000 19.240000 ;
      RECT 141.560000 18.160000 184.760000 19.240000 ;
      RECT 96.560000 18.160000 139.760000 19.240000 ;
      RECT 51.560000 18.160000 94.760000 19.240000 ;
      RECT 6.560000 18.160000 49.760000 19.240000 ;
      RECT 2.530000 18.160000 4.595000 19.240000 ;
      RECT 0.000000 18.160000 0.730000 19.240000 ;
      RECT 0.000000 16.520000 200.100000 18.160000 ;
      RECT 197.570000 15.440000 200.100000 16.520000 ;
      RECT 188.560000 15.440000 195.770000 16.520000 ;
      RECT 143.560000 15.440000 186.760000 16.520000 ;
      RECT 98.560000 15.440000 141.760000 16.520000 ;
      RECT 53.560000 15.440000 96.760000 16.520000 ;
      RECT 8.560000 15.440000 51.760000 16.520000 ;
      RECT 4.330000 15.440000 6.760000 16.520000 ;
      RECT 0.000000 15.440000 2.530000 16.520000 ;
      RECT 0.000000 13.800000 200.100000 15.440000 ;
      RECT 199.370000 12.720000 200.100000 13.800000 ;
      RECT 186.560000 12.720000 197.570000 13.800000 ;
      RECT 141.560000 12.720000 184.760000 13.800000 ;
      RECT 96.560000 12.720000 139.760000 13.800000 ;
      RECT 51.560000 12.720000 94.760000 13.800000 ;
      RECT 6.560000 12.720000 49.760000 13.800000 ;
      RECT 2.530000 12.720000 4.595000 13.800000 ;
      RECT 0.000000 12.720000 0.730000 13.800000 ;
      RECT 0.000000 11.080000 200.100000 12.720000 ;
      RECT 197.570000 10.000000 200.100000 11.080000 ;
      RECT 188.560000 10.000000 195.770000 11.080000 ;
      RECT 143.560000 10.000000 186.760000 11.080000 ;
      RECT 98.560000 10.000000 141.760000 11.080000 ;
      RECT 53.560000 10.000000 96.760000 11.080000 ;
      RECT 8.560000 10.000000 51.760000 11.080000 ;
      RECT 4.330000 10.000000 6.760000 11.080000 ;
      RECT 0.000000 10.000000 2.530000 11.080000 ;
      RECT 0.000000 8.360000 200.100000 10.000000 ;
      RECT 199.370000 7.280000 200.100000 8.360000 ;
      RECT 186.560000 7.280000 197.570000 8.360000 ;
      RECT 141.560000 7.280000 184.760000 8.360000 ;
      RECT 96.560000 7.280000 139.760000 8.360000 ;
      RECT 51.560000 7.280000 94.760000 8.360000 ;
      RECT 6.560000 7.280000 49.760000 8.360000 ;
      RECT 2.530000 7.280000 4.595000 8.360000 ;
      RECT 0.000000 7.280000 0.730000 8.360000 ;
      RECT 0.000000 5.640000 200.100000 7.280000 ;
      RECT 197.570000 4.560000 200.100000 5.640000 ;
      RECT 188.560000 4.560000 195.770000 5.640000 ;
      RECT 143.560000 4.560000 186.760000 5.640000 ;
      RECT 98.560000 4.560000 141.760000 5.640000 ;
      RECT 53.560000 4.560000 96.760000 5.640000 ;
      RECT 8.560000 4.560000 51.760000 5.640000 ;
      RECT 4.330000 4.560000 6.760000 5.640000 ;
      RECT 0.000000 4.560000 2.530000 5.640000 ;
      RECT 0.000000 4.350000 200.100000 4.560000 ;
      RECT 0.000000 0.000000 200.100000 0.750000 ;
    LAYER met4 ;
      RECT 4.330000 29.000000 195.770000 30.260000 ;
      RECT 186.560000 27.200000 195.770000 29.000000 ;
      RECT 141.560000 27.200000 184.760000 29.000000 ;
      RECT 96.560000 27.200000 139.760000 29.000000 ;
      RECT 51.560000 27.200000 94.760000 29.000000 ;
      RECT 6.560000 27.200000 49.760000 29.000000 ;
      RECT 4.330000 24.680000 4.760000 29.000000 ;
      RECT 4.330000 23.600000 4.595000 24.680000 ;
      RECT 4.330000 19.240000 4.760000 23.600000 ;
      RECT 4.330000 18.160000 4.595000 19.240000 ;
      RECT 4.330000 13.800000 4.760000 18.160000 ;
      RECT 4.330000 12.720000 4.595000 13.800000 ;
      RECT 4.330000 8.360000 4.760000 12.720000 ;
      RECT 4.330000 7.280000 4.595000 8.360000 ;
      RECT 188.560000 2.550000 195.770000 27.200000 ;
      RECT 186.560000 2.550000 186.760000 27.200000 ;
      RECT 143.560000 2.550000 184.760000 27.200000 ;
      RECT 141.560000 2.550000 141.760000 27.200000 ;
      RECT 98.560000 2.550000 139.760000 27.200000 ;
      RECT 96.560000 2.550000 96.760000 27.200000 ;
      RECT 53.560000 2.550000 94.760000 27.200000 ;
      RECT 51.560000 2.550000 51.760000 27.200000 ;
      RECT 8.560000 2.550000 49.760000 27.200000 ;
      RECT 6.560000 2.550000 6.760000 27.200000 ;
      RECT 186.560000 0.750000 195.770000 2.550000 ;
      RECT 141.560000 0.750000 184.760000 2.550000 ;
      RECT 96.560000 0.750000 139.760000 2.550000 ;
      RECT 51.560000 0.750000 94.760000 2.550000 ;
      RECT 6.560000 0.750000 49.760000 2.550000 ;
      RECT 4.330000 0.750000 4.760000 7.280000 ;
      RECT 199.370000 0.000000 200.100000 30.260000 ;
      RECT 4.330000 0.000000 195.770000 0.750000 ;
      RECT 0.000000 0.000000 0.730000 30.260000 ;
  END
END N_term_single

END LIBRARY
