##
## LEF for PtnCells ;
## created by Innovus v19.11-s128_1 on Thu Nov 25 18:57:09 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO W_IO
  CLASS BLOCK ;
  SIZE 80.040000 BY 200.260000 ;
  FOREIGN W_IO 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 80.720000 80.040000 81.100000 ;
    END
  END E1BEG[3]
  PIN E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.0224 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.448 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 79.500000 80.040000 79.880000 ;
    END
  END E1BEG[2]
  PIN E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 77.670000 80.040000 78.050000 ;
    END
  END E1BEG[1]
  PIN E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.4384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 76.450000 80.040000 76.830000 ;
    END
  END E1BEG[0]
  PIN E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 92.920000 80.040000 93.300000 ;
    END
  END E2BEG[7]
  PIN E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.9244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.592 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 91.090000 80.040000 91.470000 ;
    END
  END E2BEG[6]
  PIN E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 89.870000 80.040000 90.250000 ;
    END
  END E2BEG[5]
  PIN E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 88.040000 80.040000 88.420000 ;
    END
  END E2BEG[4]
  PIN E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 86.820000 80.040000 87.200000 ;
    END
  END E2BEG[3]
  PIN E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.1044 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.552 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 84.990000 80.040000 85.370000 ;
    END
  END E2BEG[2]
  PIN E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 83.770000 80.040000 84.150000 ;
    END
  END E2BEG[1]
  PIN E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 81.940000 80.040000 82.320000 ;
    END
  END E2BEG[0]
  PIN E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 104.510000 80.040000 104.890000 ;
    END
  END E2BEGb[7]
  PIN E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 103.290000 80.040000 103.670000 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 101.460000 80.040000 101.840000 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 100.240000 80.040000 100.620000 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 98.410000 80.040000 98.790000 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.6694 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 94.232 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 97.190000 80.040000 97.570000 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 95.360000 80.040000 95.740000 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 94.140000 80.040000 94.520000 ;
    END
  END E2BEGb[0]
  PIN EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 128.300000 80.040000 128.680000 ;
    END
  END EE4BEG[15]
  PIN EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.3308 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.568 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 127.080000 80.040000 127.460000 ;
    END
  END EE4BEG[14]
  PIN EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 125.250000 80.040000 125.630000 ;
    END
  END EE4BEG[13]
  PIN EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.2164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.816 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 124.030000 80.040000 124.410000 ;
    END
  END EE4BEG[12]
  PIN EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 122.200000 80.040000 122.580000 ;
    END
  END EE4BEG[11]
  PIN EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.0934 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.16 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 120.980000 80.040000 121.360000 ;
    END
  END EE4BEG[10]
  PIN EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 119.150000 80.040000 119.530000 ;
    END
  END EE4BEG[9]
  PIN EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 117.930000 80.040000 118.310000 ;
    END
  END EE4BEG[8]
  PIN EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.5194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.432 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 116.710000 80.040000 117.090000 ;
    END
  END EE4BEG[7]
  PIN EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.3924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.088 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 114.880000 80.040000 115.260000 ;
    END
  END EE4BEG[6]
  PIN EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 113.660000 80.040000 114.040000 ;
    END
  END EE4BEG[5]
  PIN EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.0584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 111.830000 80.040000 112.210000 ;
    END
  END EE4BEG[4]
  PIN EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.9594 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.112 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 110.610000 80.040000 110.990000 ;
    END
  END EE4BEG[3]
  PIN EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.3862 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.192 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 108.780000 80.040000 109.160000 ;
    END
  END EE4BEG[2]
  PIN EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 107.560000 80.040000 107.940000 ;
    END
  END EE4BEG[1]
  PIN EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 105.730000 80.040000 106.110000 ;
    END
  END EE4BEG[0]
  PIN E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 145.990000 80.040000 146.370000 ;
    END
  END E6BEG[11]
  PIN E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.4764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.536 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 144.770000 80.040000 145.150000 ;
    END
  END E6BEG[10]
  PIN E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 143.550000 80.040000 143.930000 ;
    END
  END E6BEG[9]
  PIN E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.9224 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.248 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 141.720000 80.040000 142.100000 ;
    END
  END E6BEG[8]
  PIN E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 140.500000 80.040000 140.880000 ;
    END
  END E6BEG[7]
  PIN E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.9388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.144 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 138.670000 80.040000 139.050000 ;
    END
  END E6BEG[6]
  PIN E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.3684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.96 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 137.450000 80.040000 137.830000 ;
    END
  END E6BEG[5]
  PIN E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 135.620000 80.040000 136.000000 ;
    END
  END E6BEG[4]
  PIN E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 134.400000 80.040000 134.780000 ;
    END
  END E6BEG[3]
  PIN E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 132.570000 80.040000 132.950000 ;
    END
  END E6BEG[2]
  PIN E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 131.350000 80.040000 131.730000 ;
    END
  END E6BEG[1]
  PIN E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 130.130000 80.040000 130.510000 ;
    END
  END E6BEG[0]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.9412 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.152 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8787 LAYER met3  ;
    ANTENNAMAXAREACAR 44.2498 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 212.659 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.550615 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 9.350000 80.040000 9.730000 ;
    END
  END W1END[3]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.7408 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.088 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8787 LAYER met3  ;
    ANTENNAMAXAREACAR 36.2681 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 163.762 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 7.520000 80.040000 7.900000 ;
    END
  END W1END[2]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.7224 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.648 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met3  ;
    ANTENNAMAXAREACAR 44.4845 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 214.494 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.621955 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.936 LAYER met4  ;
    ANTENNAGATEAREA 0.8787 LAYER met4  ;
    ANTENNAMAXAREACAR 46.0776 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 223.526 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 6.300000 80.040000 6.680000 ;
    END
  END W1END[1]
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.104 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 17.8242 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 71.9036 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.3237 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 162.192 LAYER met4  ;
    ANTENNAGATEAREA 0.8787 LAYER met4  ;
    ANTENNAMAXAREACAR 52.334 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 256.485 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 5.080000 80.040000 5.460000 ;
    END
  END W1END[0]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.3924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.088 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5477 LAYER met3  ;
    ANTENNAMAXAREACAR 47.3066 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 228.811 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.773644 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 20.940000 80.040000 21.320000 ;
    END
  END W2MID[7]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.4342 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met3  ;
    ANTENNAMAXAREACAR 33.6968 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 153.168 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.411019 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 19.720000 80.040000 20.100000 ;
    END
  END W2MID[6]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.436 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.792 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 28.8392 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 127.467 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.482697 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.2558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.168 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 34.7397 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 159.318 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.490985 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 17.890000 80.040000 18.270000 ;
    END
  END W2MID[5]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met3  ;
    ANTENNAMAXAREACAR 25.8056 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 110.752 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.355799 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 16.670000 80.040000 17.050000 ;
    END
  END W2MID[4]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.3434 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.16 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met3  ;
    ANTENNAMAXAREACAR 31.5387 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 148.371 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.497308 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 15.450000 80.040000 15.830000 ;
    END
  END W2MID[3]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4624 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met3  ;
    ANTENNAMAXAREACAR 27.851 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 120.331 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.497308 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 13.620000 80.040000 14.000000 ;
    END
  END W2MID[2]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met3  ;
    ANTENNAMAXAREACAR 31.2345 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 137.44 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.497308 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 12.400000 80.040000 12.780000 ;
    END
  END W2MID[1]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.3704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.104 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 35.4276 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 166.97 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.525393 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.9378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.472 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 42.2441 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 210.902 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.637736 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 10.570000 80.040000 10.950000 ;
    END
  END W2MID[0]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.2132 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.936 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0707 LAYER met3  ;
    ANTENNAMAXAREACAR 36.0551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 168.009 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 33.140000 80.040000 33.520000 ;
    END
  END W2END[7]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.3311 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.56 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met3  ;
    ANTENNAMAXAREACAR 77.3686 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 381.267 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 31.310000 80.040000 31.690000 ;
    END
  END W2END[6]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.8263 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.064 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met3  ;
    ANTENNAMAXAREACAR 35.3148 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 173.642 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.515094 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 30.090000 80.040000 30.470000 ;
    END
  END W2END[5]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.072 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met3  ;
    ANTENNAMAXAREACAR 30.5771 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 134.218 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.352074 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 28.870000 80.040000 29.250000 ;
    END
  END W2END[4]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.1949 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 119.304 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met3  ;
    ANTENNAMAXAREACAR 39.3281 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 197.614 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 27.040000 80.040000 27.420000 ;
    END
  END W2END[3]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.4191 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.696 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met3  ;
    ANTENNAMAXAREACAR 26.9854 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 122.231 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 25.820000 80.040000 26.200000 ;
    END
  END W2END[2]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met3  ;
    ANTENNAMAXAREACAR 27.0875 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 116.465 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.355799 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 23.990000 80.040000 24.370000 ;
    END
  END W2END[1]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.426 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met3  ;
    ANTENNAMAXAREACAR 40.9567 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 199.207 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 22.770000 80.040000 23.150000 ;
    END
  END W2END[0]
  PIN WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.2922 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 24.4798 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 106.323 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 56.930000 80.040000 57.310000 ;
    END
  END WW4END[15]
  PIN WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.9884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 16.915 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 66.6132 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367145 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 55.100000 80.040000 55.480000 ;
    END
  END WW4END[14]
  PIN WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 16.4444 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 74.4971 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367145 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 53.880000 80.040000 54.260000 ;
    END
  END WW4END[13]
  PIN WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 13.5729 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 50.4684 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.525393 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.7568 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 57.84 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 25.3715 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 113.91 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 52.660000 80.040000 53.040000 ;
    END
  END WW4END[12]
  PIN WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.5984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.52 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 29.7621 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 132.511 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367145 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 50.830000 80.040000 51.210000 ;
    END
  END WW4END[11]
  PIN WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.4942 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 31.2363 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 141.05 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 49.610000 80.040000 49.990000 ;
    END
  END WW4END[10]
  PIN WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.0181 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.224 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 51.3943 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 255.743 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 47.780000 80.040000 48.160000 ;
    END
  END WW4END[9]
  PIN WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.572 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.32 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 35.6576 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 161.562 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 46.560000 80.040000 46.940000 ;
    END
  END WW4END[8]
  PIN WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.8744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.992 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 25.9781 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 124.312 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.508654 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 44.730000 80.040000 45.110000 ;
    END
  END WW4END[7]
  PIN WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 17.3798 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 68.1934 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.508654 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 43.510000 80.040000 43.890000 ;
    END
  END WW4END[6]
  PIN WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.6765 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.928 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 42.8111 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 208.673 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.0225 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 97.056 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 62.5792 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 315.129 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 42.290000 80.040000 42.670000 ;
    END
  END WW4END[5]
  PIN WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 20.4873 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 83.6178 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367145 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 40.460000 80.040000 40.840000 ;
    END
  END WW4END[4]
  PIN WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.9012 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.272 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 30.8429 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 147.824 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.458019 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 39.240000 80.040000 39.620000 ;
    END
  END WW4END[3]
  PIN WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 23.717 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 100.283 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.508654 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 37.410000 80.040000 37.790000 ;
    END
  END WW4END[2]
  PIN WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.8895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.064 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 37.1799 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 178.473 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.7666 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 79.696 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 53.3767 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 265.887 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 36.190000 80.040000 36.570000 ;
    END
  END WW4END[1]
  PIN WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 28.2509 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 133.33 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367145 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 34.360000 80.040000 34.740000 ;
    END
  END WW4END[0]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7866 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.0858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.928 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 32.2185 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 162.634 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.411019 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 74.620000 80.040000 75.000000 ;
    END
  END W6END[11]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.9128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.672 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0707 LAYER met3  ;
    ANTENNAMAXAREACAR 15.6999 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 73.1544 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 73.400000 80.040000 73.780000 ;
    END
  END W6END[10]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.558 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.432 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 38.1242 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 178.164 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 71.570000 80.040000 71.950000 ;
    END
  END W6END[9]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1846 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.976 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.3668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 55.76 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0707 LAYER met4  ;
    ANTENNAMAXAREACAR 29.8352 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 146.898 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.612202 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 70.350000 80.040000 70.730000 ;
    END
  END W6END[8]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.344 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.104 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met3  ;
    ANTENNAMAXAREACAR 32.6765 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 149.06 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 68.520000 80.040000 68.900000 ;
    END
  END W6END[7]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met3  ;
    ANTENNAMAXAREACAR 29.0092 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 138.989 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.493584 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 67.300000 80.040000 67.680000 ;
    END
  END W6END[6]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3726 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.5848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.256 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 32.5589 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 162.893 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.522388 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 66.080000 80.040000 66.460000 ;
    END
  END W6END[5]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met3  ;
    ANTENNAMAXAREACAR 32.2984 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 155.357 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.493584 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 64.250000 80.040000 64.630000 ;
    END
  END W6END[4]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.9659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met3  ;
    ANTENNAMAXAREACAR 40.1763 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 197.815 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 63.030000 80.040000 63.410000 ;
    END
  END W6END[3]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met3  ;
    ANTENNAMAXAREACAR 23.0253 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 107.999 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.497308 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 61.200000 80.040000 61.580000 ;
    END
  END W6END[2]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.9444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.032 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met3  ;
    ANTENNAMAXAREACAR 36.3494 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 178.152 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.493584 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 59.980000 80.040000 60.360000 ;
    END
  END W6END[1]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.6529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.472 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 15.4198 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 60.5163 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.458019 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.2688 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 49.904 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 42.8348 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 214.182 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.695388 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 58.150000 80.040000 58.530000 ;
    END
  END W6END[0]
  PIN A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.1964 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.376 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 42.290000 0.700000 42.670000 ;
    END
  END A_I_top
  PIN A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 38.630000 0.700000 39.010000 ;
    END
  END A_T_top
  PIN A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3751 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.128 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.4817 LAYER met3  ;
    ANTENNAMAXAREACAR 30.21 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 146.075 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.729187 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 34.360000 0.700000 34.740000 ;
    END
  END A_O_top
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9492 LAYER met3  ;
    ANTENNAMAXAREACAR 16.2608 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 67.167 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.365411 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 0.000000 5.480000 0.700000 ;
    END
  END UserCLK
  PIN B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 13.010000 0.700000 13.390000 ;
    END
  END B_I_top
  PIN B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 8.740000 0.700000 9.120000 ;
    END
  END B_T_top
  PIN B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.4682 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 94.096 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8457 LAYER met3  ;
    ANTENNAMAXAREACAR 42.6692 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 211.331 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.914508 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.1708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.048 LAYER met4  ;
    ANTENNAGATEAREA 1.4817 LAYER met4  ;
    ANTENNAMAXAREACAR 48.1837 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 241.059 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.914508 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 5.080000 0.700000 5.460000 ;
    END
  END B_O_top
  PIN A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 46.560000 0.700000 46.940000 ;
    END
  END A_config_C_bit0
  PIN A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 50.830000 0.700000 51.210000 ;
    END
  END A_config_C_bit1
  PIN A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.6784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 55.100000 0.700000 55.480000 ;
    END
  END A_config_C_bit2
  PIN A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 59.370000 0.700000 59.750000 ;
    END
  END A_config_C_bit3
  PIN B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 17.280000 0.700000 17.660000 ;
    END
  END B_config_C_bit0
  PIN B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 21.550000 0.700000 21.930000 ;
    END
  END B_config_C_bit1
  PIN B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 25.820000 0.700000 26.200000 ;
    END
  END B_config_C_bit2
  PIN B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 30.090000 0.700000 30.470000 ;
    END
  END B_config_C_bit3
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3488 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.734 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 199.560000 5.480000 200.260000 ;
    END
  END UserCLKo
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6392 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.688 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met3  ;
    ANTENNAMAXAREACAR 63.4706 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 318.582 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 194.180000 0.700000 194.560000 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.368 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met3  ;
    ANTENNAMAXAREACAR 32.6655 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 159.852 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.371318 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 189.910000 0.700000 190.290000 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.4391 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 168.616 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met3  ;
    ANTENNAMAXAREACAR 83.6414 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 426.63 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.632495 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 185.640000 0.700000 186.020000 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4518 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.68 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3555 LAYER met3  ;
    ANTENNAMAXAREACAR 97.8697 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.895724 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.9777 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 101.68 LAYER met4  ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 120.666 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 613.218 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.895724 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 181.370000 0.700000 181.750000 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.0942 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.776 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5145 LAYER met3  ;
    ANTENNAMAXAREACAR 61.1226 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 308.21 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.794098 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.5628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.472 LAYER met4  ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 76.213 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 389.257 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.794098 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 177.100000 0.700000 177.480000 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.94935 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.936 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 56.1626 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 282.237 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.986768 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 36.4347 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 194.784 LAYER met4  ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 99.928 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 516.211 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.986768 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 172.830000 0.700000 173.210000 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.0392 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.7552 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 176.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 71.4838 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 372.404 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 168.560000 0.700000 168.940000 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.6817 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.248 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met3  ;
    ANTENNAMAXAREACAR 42.3078 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 211.055 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.449057 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 164.290000 0.700000 164.670000 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.536 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 80.3644 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 424.356 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 25.2618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 135.2 LAYER met4  ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 110.709 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 586.759 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 160.020000 0.700000 160.400000 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1393 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.688 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 30.9888 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 159.865 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.872265 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.8238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 148.864 LAYER met4  ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 64.4108 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 338.681 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.872265 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 155.750000 0.700000 156.130000 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.152 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3555 LAYER met3  ;
    ANTENNAMAXAREACAR 65.0425 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 329.766 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.660823 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 25.4688 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 136.304 LAYER met4  ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 95.6357 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 493.494 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.660823 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 152.090000 0.700000 152.470000 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.936 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 86.888 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 445.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.4971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 179.112 LAYER met4  ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 127.125 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 661.094 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 147.820000 0.700000 148.200000 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5089 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.656 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3555 LAYER met3  ;
    ANTENNAMAXAREACAR 59.5738 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 296.284 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.802333 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.9577 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 160.24 LAYER met4  ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 95.559 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 488.765 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 143.550000 0.700000 143.930000 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.52 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3555 LAYER met3  ;
    ANTENNAMAXAREACAR 68.5524 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 346.325 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.660823 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.6108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.728 LAYER met4  ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 83.7005 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 427.68 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.660823 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 139.280000 0.700000 139.660000 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5085 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.032 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 64.4868 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 327.421 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.6319 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 64.384 LAYER met4  ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 78.459 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 404.76 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 135.010000 0.700000 135.390000 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.6972 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.2416 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 60.896 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 81.7833 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 426.504 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700629 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 130.740000 0.700000 131.120000 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.104 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met3  ;
    ANTENNAMAXAREACAR 60.5427 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 298.682 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.512828 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 126.470000 0.700000 126.850000 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met3  ;
    ANTENNAMAXAREACAR 42.0721 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 206.476 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.857862 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.6438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.904 LAYER met4  ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 46.4491 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 230.385 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.857862 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 122.200000 0.700000 122.580000 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.7442 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met3  ;
    ANTENNAMAXAREACAR 64.9631 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 331.536 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 117.930000 0.700000 118.310000 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.8663 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 106.424 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met3  ;
    ANTENNAMAXAREACAR 48.0072 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 246.045 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 114.270000 0.700000 114.650000 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.0661 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.96 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met3  ;
    ANTENNAMAXAREACAR 47.6787 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 241.278 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 110.000000 0.700000 110.380000 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1089 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.056 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met3  ;
    ANTENNAMAXAREACAR 43.07 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 211.219 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.524171 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 105.730000 0.700000 106.110000 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.936 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met3  ;
    ANTENNAMAXAREACAR 60.0305 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 297.139 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.524171 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 101.460000 0.700000 101.840000 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.9422 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.304 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met3  ;
    ANTENNAMAXAREACAR 43.9195 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 223.127 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 97.190000 0.700000 97.570000 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.352 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met3  ;
    ANTENNAMAXAREACAR 38.071 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 187.198 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.665681 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 92.920000 0.700000 93.300000 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4697 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.784 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met3  ;
    ANTENNAMAXAREACAR 22.8199 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 111.284 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 88.650000 0.700000 89.030000 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6417 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.368 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met3  ;
    ANTENNAMAXAREACAR 58.5691 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 288.995 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 84.380000 0.700000 84.760000 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.9605 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.776 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 82.8679 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 434.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.4726 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.128 LAYER met4  ;
    ANTENNAGATEAREA 0.6735 LAYER met4  ;
    ANTENNAMAXAREACAR 95.4479 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 503.298 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 80.110000 0.700000 80.490000 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.8491 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.136 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met3  ;
    ANTENNAMAXAREACAR 50.9691 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 257.091 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 76.450000 0.700000 76.830000 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6972 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.664 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met3  ;
    ANTENNAMAXAREACAR 49.4532 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 245.289 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.620271 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 72.180000 0.700000 72.560000 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.3645 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 98.88 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met4  ;
    ANTENNAMAXAREACAR 59.1943 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 304.33 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.689815 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 67.910000 0.700000 68.290000 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.3162 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 92.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.5223 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 132.192 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met4  ;
    ANTENNAMAXAREACAR 61.1707 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 318.803 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 63.640000 0.700000 64.020000 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.6324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.368 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 194.180000 80.040000 194.560000 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 192.350000 80.040000 192.730000 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.0584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 191.130000 80.040000 191.510000 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 189.300000 80.040000 189.680000 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.0584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 188.080000 80.040000 188.460000 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.9544 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.752 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 186.250000 80.040000 186.630000 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 185.030000 80.040000 185.410000 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.1264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.336 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 183.200000 80.040000 183.580000 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 181.980000 80.040000 182.360000 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.9904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.944 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 180.760000 80.040000 181.140000 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 178.930000 80.040000 179.310000 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.6104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.584 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 177.710000 80.040000 178.090000 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 175.880000 80.040000 176.260000 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.2664 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.416 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 174.660000 80.040000 175.040000 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.3344 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.112 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 172.830000 80.040000 173.210000 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.6784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 171.610000 80.040000 171.990000 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 169.780000 80.040000 170.160000 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 168.560000 80.040000 168.940000 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.6784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 167.340000 80.040000 167.720000 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 165.510000 80.040000 165.890000 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.8524 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.208 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 164.290000 80.040000 164.670000 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 162.460000 80.040000 162.840000 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.6104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.584 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 161.240000 80.040000 161.620000 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 159.410000 80.040000 159.790000 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.1304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.024 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 158.190000 80.040000 158.570000 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.3384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.8 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 156.360000 80.040000 156.740000 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.0224 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.256 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 155.140000 80.040000 155.520000 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 153.920000 80.040000 154.300000 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.5414 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.216 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 152.090000 80.040000 152.470000 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.2324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.568 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 150.870000 80.040000 151.250000 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 149.040000 80.040000 149.420000 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 79.340000 147.820000 80.040000 148.200000 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.9505 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 119.592 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.5588 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.784 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 31.1858 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 165.109 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 74.560000 0.000000 74.940000 0.700000 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7809 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.7435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.7397 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 201.744 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 92.8132 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 471.824 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 70.880000 0.000000 71.260000 0.700000 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.9047 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 266.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 101.974 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 524.388 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 67.200000 0.000000 67.580000 0.700000 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.1698 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 193.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 115.331 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 595.836 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.732074 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 63.980000 0.000000 64.360000 0.700000 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6817 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.6477 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 275.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 99.4768 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 508.415 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 60.300000 0.000000 60.680000 0.700000 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7175 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.1848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 241.456 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 110.66 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 578.77 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.732074 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 57.080000 0.000000 57.460000 0.700000 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8773 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.2255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.1467 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 241.248 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 90.8838 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 462.792 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 53.400000 0.000000 53.780000 0.700000 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9737 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.7217 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 265.648 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 99.9753 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 515.281 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 50.180000 0.000000 50.560000 0.700000 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6817 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.1577 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 246.64 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 87.7181 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 448.926 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 46.500000 0.000000 46.880000 0.700000 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7175 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.8558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 234.368 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 79.3199 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 403.496 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.38832 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 43.280000 0.000000 43.660000 0.700000 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5109 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.3935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.5717 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 232.848 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 77.3619 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 394.142 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 39.600000 0.000000 39.980000 0.700000 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4255 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.9665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.5488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 222.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 73.5411 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 373.154 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.38832 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 35.920000 0.000000 36.300000 0.700000 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4503 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.0905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.9258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 197.408 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 64.8321 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 327.408 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.309463 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 32.700000 0.000000 33.080000 0.700000 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0915 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.2965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.8397 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 228.944 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 76.2549 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 387.674 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 29.020000 0.000000 29.400000 0.700000 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2795 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.2365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.0357 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 224.656 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 80.8168 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 428.046 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 25.800000 0.000000 26.180000 0.700000 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0839 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.1568 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 182.64 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 68.9461 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 348.461 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.38832 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 22.120000 0.000000 22.500000 0.700000 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.5463 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.0105 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0707 LAYER met2  ;
    ANTENNAMAXAREACAR 14.8927 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 69.2302 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.502139 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.4696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.112 LAYER met3  ;
    ANTENNAGATEAREA 3.4932 LAYER met3  ;
    ANTENNAMAXAREACAR 19.5704 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 93.0762 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.534315 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 18.900000 0.000000 19.280000 0.700000 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 30.236 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 147.868 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.7192 LAYER met2  ;
    ANTENNAMAXAREACAR 24.6572 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 117.043 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.606289 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 15.220000 0.000000 15.600000 0.700000 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 18.0334 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 88.361 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3427 LAYER met2  ;
    ANTENNAMAXAREACAR 15.9084 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 73.7868 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.498929 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.3535 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.488 LAYER met3  ;
    ANTENNAGATEAREA 5.7192 LAYER met3  ;
    ANTENNAMAXAREACAR 19.978 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 94.1194 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.619368 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 12.000000 0.000000 12.380000 0.700000 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 28.5584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 139.748 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.7652 LAYER met2  ;
    ANTENNAMAXAREACAR 31.2104 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 150.673 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.663329 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.1394 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 135.008 LAYER met3  ;
    ANTENNAGATEAREA 5.7192 LAYER met3  ;
    ANTENNAMAXAREACAR 35.606 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 174.279 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.663329 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 8.320000 0.000000 8.700000 0.700000 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9382 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.583 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 74.560000 199.560000 74.940000 200.260000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5574 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.679 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 70.880000 199.560000 71.260000 200.260000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4342 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.063 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 67.200000 199.560000 67.580000 200.260000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.129 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.537 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 63.980000 199.560000 64.360000 200.260000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.431 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 60.300000 199.560000 60.680000 200.260000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3834 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.809 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 57.080000 199.560000 57.460000 200.260000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.319 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.487 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 53.400000 199.560000 53.780000 200.260000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.971 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.747 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 50.180000 199.560000 50.560000 200.260000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8422 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.103 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 46.500000 199.560000 46.880000 200.260000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.2866 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.325 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 43.280000 199.560000 43.660000 200.260000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.6874 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.329 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 39.600000 199.560000 39.980000 200.260000 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.6198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.991 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 35.920000 199.560000 36.300000 200.260000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.3394 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.589 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 32.700000 199.560000 33.080000 200.260000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.9066 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 29.020000 199.560000 29.400000 200.260000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0354 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.069 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 25.800000 199.560000 26.180000 200.260000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.223 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.007 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 22.120000 199.560000 22.500000 200.260000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.4602 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.193 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 18.900000 199.560000 19.280000 200.260000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.5586 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.685 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 15.220000 199.560000 15.600000 200.260000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.971 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.747 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 12.000000 199.560000 12.380000 200.260000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.9066 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 8.320000 199.560000 8.700000 200.260000 ;
    END
  END FrameStrobe_O[0]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 78.840000 195.020000 80.040000 196.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 195.020000 1.200000 196.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.840000 2.850000 80.040000 4.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 1.200000 4.050000 ;
    END
    PORT
      LAYER met4 ;
        RECT 76.010000 199.060000 77.210000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 76.010000 0.000000 77.210000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 199.060000 4.030000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 0.000000 4.030000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 80.040000 4.050000 ;
        RECT 0.000000 195.020000 80.040000 196.220000 ;
        RECT 2.830000 4.860000 4.030000 5.340000 ;
        RECT 2.830000 10.300000 4.030000 10.780000 ;
        RECT 7.060000 10.300000 8.260000 10.780000 ;
        RECT 7.060000 4.860000 8.260000 5.340000 ;
        RECT 7.060000 21.180000 8.260000 21.660000 ;
        RECT 7.060000 15.740000 8.260000 16.220000 ;
        RECT 2.830000 21.180000 4.030000 21.660000 ;
        RECT 2.830000 15.740000 4.030000 16.220000 ;
        RECT 2.830000 37.500000 4.030000 37.980000 ;
        RECT 7.060000 37.500000 8.260000 37.980000 ;
        RECT 7.060000 32.060000 8.260000 32.540000 ;
        RECT 7.060000 26.620000 8.260000 27.100000 ;
        RECT 2.830000 32.060000 4.030000 32.540000 ;
        RECT 2.830000 26.620000 4.030000 27.100000 ;
        RECT 7.060000 48.380000 8.260000 48.860000 ;
        RECT 7.060000 42.940000 8.260000 43.420000 ;
        RECT 2.830000 48.380000 4.030000 48.860000 ;
        RECT 2.830000 42.940000 4.030000 43.420000 ;
        RECT 7.060000 53.820000 8.260000 54.300000 ;
        RECT 7.060000 59.260000 8.260000 59.740000 ;
        RECT 2.830000 59.260000 4.030000 59.740000 ;
        RECT 2.830000 53.820000 4.030000 54.300000 ;
        RECT 7.060000 64.700000 8.260000 65.180000 ;
        RECT 7.060000 70.140000 8.260000 70.620000 ;
        RECT 2.830000 70.140000 4.030000 70.620000 ;
        RECT 2.830000 64.700000 4.030000 65.180000 ;
        RECT 7.060000 81.020000 8.260000 81.500000 ;
        RECT 2.830000 81.020000 4.030000 81.500000 ;
        RECT 2.830000 75.580000 4.030000 76.060000 ;
        RECT 7.060000 75.580000 8.260000 76.060000 ;
        RECT 2.830000 86.460000 4.030000 86.940000 ;
        RECT 7.060000 86.460000 8.260000 86.940000 ;
        RECT 7.060000 91.900000 8.260000 92.380000 ;
        RECT 7.060000 97.340000 8.260000 97.820000 ;
        RECT 2.830000 97.340000 4.030000 97.820000 ;
        RECT 2.830000 91.900000 4.030000 92.380000 ;
        RECT 52.060000 21.180000 53.260000 21.660000 ;
        RECT 52.060000 4.860000 53.260000 5.340000 ;
        RECT 52.060000 10.300000 53.260000 10.780000 ;
        RECT 52.060000 15.740000 53.260000 16.220000 ;
        RECT 76.010000 10.300000 77.210000 10.780000 ;
        RECT 76.010000 4.860000 77.210000 5.340000 ;
        RECT 76.010000 21.180000 77.210000 21.660000 ;
        RECT 76.010000 15.740000 77.210000 16.220000 ;
        RECT 52.060000 48.380000 53.260000 48.860000 ;
        RECT 52.060000 42.940000 53.260000 43.420000 ;
        RECT 52.060000 37.500000 53.260000 37.980000 ;
        RECT 52.060000 32.060000 53.260000 32.540000 ;
        RECT 52.060000 26.620000 53.260000 27.100000 ;
        RECT 76.010000 37.500000 77.210000 37.980000 ;
        RECT 76.010000 32.060000 77.210000 32.540000 ;
        RECT 76.010000 26.620000 77.210000 27.100000 ;
        RECT 76.010000 48.380000 77.210000 48.860000 ;
        RECT 76.010000 42.940000 77.210000 43.420000 ;
        RECT 52.060000 53.820000 53.260000 54.300000 ;
        RECT 52.060000 59.260000 53.260000 59.740000 ;
        RECT 52.060000 64.700000 53.260000 65.180000 ;
        RECT 52.060000 70.140000 53.260000 70.620000 ;
        RECT 76.010000 59.260000 77.210000 59.740000 ;
        RECT 76.010000 53.820000 77.210000 54.300000 ;
        RECT 76.010000 70.140000 77.210000 70.620000 ;
        RECT 76.010000 64.700000 77.210000 65.180000 ;
        RECT 52.060000 75.580000 53.260000 76.060000 ;
        RECT 52.060000 81.020000 53.260000 81.500000 ;
        RECT 52.060000 86.460000 53.260000 86.940000 ;
        RECT 52.060000 91.900000 53.260000 92.380000 ;
        RECT 52.060000 97.340000 53.260000 97.820000 ;
        RECT 76.010000 86.460000 77.210000 86.940000 ;
        RECT 76.010000 81.020000 77.210000 81.500000 ;
        RECT 76.010000 75.580000 77.210000 76.060000 ;
        RECT 76.010000 97.340000 77.210000 97.820000 ;
        RECT 76.010000 91.900000 77.210000 92.380000 ;
        RECT 7.060000 102.780000 8.260000 103.260000 ;
        RECT 7.060000 108.220000 8.260000 108.700000 ;
        RECT 2.830000 108.220000 4.030000 108.700000 ;
        RECT 2.830000 102.780000 4.030000 103.260000 ;
        RECT 2.830000 113.660000 4.030000 114.140000 ;
        RECT 7.060000 113.660000 8.260000 114.140000 ;
        RECT 2.830000 119.100000 4.030000 119.580000 ;
        RECT 2.830000 124.540000 4.030000 125.020000 ;
        RECT 7.060000 119.100000 8.260000 119.580000 ;
        RECT 7.060000 124.540000 8.260000 125.020000 ;
        RECT 7.060000 135.420000 8.260000 135.900000 ;
        RECT 7.060000 129.980000 8.260000 130.460000 ;
        RECT 2.830000 135.420000 4.030000 135.900000 ;
        RECT 2.830000 129.980000 4.030000 130.460000 ;
        RECT 7.060000 146.300000 8.260000 146.780000 ;
        RECT 7.060000 140.860000 8.260000 141.340000 ;
        RECT 2.830000 146.300000 4.030000 146.780000 ;
        RECT 2.830000 140.860000 4.030000 141.340000 ;
        RECT 2.830000 162.620000 4.030000 163.100000 ;
        RECT 7.060000 162.620000 8.260000 163.100000 ;
        RECT 7.060000 151.740000 8.260000 152.220000 ;
        RECT 7.060000 157.180000 8.260000 157.660000 ;
        RECT 2.830000 157.180000 4.030000 157.660000 ;
        RECT 2.830000 151.740000 4.030000 152.220000 ;
        RECT 7.060000 168.060000 8.260000 168.540000 ;
        RECT 7.060000 173.500000 8.260000 173.980000 ;
        RECT 2.830000 173.500000 4.030000 173.980000 ;
        RECT 2.830000 168.060000 4.030000 168.540000 ;
        RECT 2.830000 184.380000 4.030000 184.860000 ;
        RECT 7.060000 178.940000 8.260000 179.420000 ;
        RECT 7.060000 184.380000 8.260000 184.860000 ;
        RECT 2.830000 178.940000 4.030000 179.420000 ;
        RECT 2.830000 189.820000 4.030000 190.300000 ;
        RECT 7.060000 189.820000 8.260000 190.300000 ;
        RECT 52.060000 124.540000 53.260000 125.020000 ;
        RECT 52.060000 119.100000 53.260000 119.580000 ;
        RECT 52.060000 102.780000 53.260000 103.260000 ;
        RECT 52.060000 108.220000 53.260000 108.700000 ;
        RECT 52.060000 113.660000 53.260000 114.140000 ;
        RECT 76.010000 108.220000 77.210000 108.700000 ;
        RECT 76.010000 102.780000 77.210000 103.260000 ;
        RECT 76.010000 124.540000 77.210000 125.020000 ;
        RECT 76.010000 119.100000 77.210000 119.580000 ;
        RECT 76.010000 113.660000 77.210000 114.140000 ;
        RECT 52.060000 146.300000 53.260000 146.780000 ;
        RECT 52.060000 140.860000 53.260000 141.340000 ;
        RECT 52.060000 135.420000 53.260000 135.900000 ;
        RECT 52.060000 129.980000 53.260000 130.460000 ;
        RECT 76.010000 135.420000 77.210000 135.900000 ;
        RECT 76.010000 129.980000 77.210000 130.460000 ;
        RECT 76.010000 146.300000 77.210000 146.780000 ;
        RECT 76.010000 140.860000 77.210000 141.340000 ;
        RECT 52.060000 151.740000 53.260000 152.220000 ;
        RECT 52.060000 157.180000 53.260000 157.660000 ;
        RECT 52.060000 162.620000 53.260000 163.100000 ;
        RECT 52.060000 168.060000 53.260000 168.540000 ;
        RECT 52.060000 173.500000 53.260000 173.980000 ;
        RECT 76.010000 162.620000 77.210000 163.100000 ;
        RECT 76.010000 157.180000 77.210000 157.660000 ;
        RECT 76.010000 151.740000 77.210000 152.220000 ;
        RECT 76.010000 173.500000 77.210000 173.980000 ;
        RECT 76.010000 168.060000 77.210000 168.540000 ;
        RECT 52.060000 178.940000 53.260000 179.420000 ;
        RECT 52.060000 184.380000 53.260000 184.860000 ;
        RECT 52.060000 189.820000 53.260000 190.300000 ;
        RECT 76.010000 184.380000 77.210000 184.860000 ;
        RECT 76.010000 178.940000 77.210000 179.420000 ;
        RECT 76.010000 189.820000 77.210000 190.300000 ;
      LAYER met4 ;
        RECT 52.060000 2.850000 53.260000 196.220000 ;
        RECT 7.060000 2.850000 8.260000 196.220000 ;
        RECT 76.010000 0.000000 77.210000 200.260000 ;
        RECT 2.830000 0.000000 4.030000 200.260000 ;
    END
# end of P/G power stripe data as pin

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 78.840000 196.820000 80.040000 198.020000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 196.820000 1.200000 198.020000 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.840000 1.050000 80.040000 2.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 1.200000 2.250000 ;
    END
    PORT
      LAYER met4 ;
        RECT 77.810000 199.060000 79.010000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 77.810000 0.000000 79.010000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 199.060000 2.230000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 0.000000 2.230000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 80.040000 2.250000 ;
        RECT 0.000000 196.820000 80.040000 198.020000 ;
        RECT 77.810000 100.060000 79.010000 100.540000 ;
        RECT 4.895000 100.060000 6.260000 100.540000 ;
        RECT 1.030000 100.060000 2.230000 100.540000 ;
        RECT 50.060000 100.060000 51.260000 100.540000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 1.030000 7.580000 2.230000 8.060000 ;
        RECT 1.030000 23.900000 2.230000 24.380000 ;
        RECT 1.030000 18.460000 2.230000 18.940000 ;
        RECT 1.030000 13.020000 2.230000 13.500000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 1.030000 29.340000 2.230000 29.820000 ;
        RECT 1.030000 34.780000 2.230000 35.260000 ;
        RECT 4.895000 29.340000 6.260000 29.820000 ;
        RECT 4.895000 34.780000 6.260000 35.260000 ;
        RECT 1.030000 40.220000 2.230000 40.700000 ;
        RECT 1.030000 45.660000 2.230000 46.140000 ;
        RECT 4.895000 40.220000 6.260000 40.700000 ;
        RECT 4.895000 45.660000 6.260000 46.140000 ;
        RECT 1.030000 61.980000 2.230000 62.460000 ;
        RECT 1.030000 56.540000 2.230000 57.020000 ;
        RECT 1.030000 51.100000 2.230000 51.580000 ;
        RECT 4.895000 61.980000 6.260000 62.460000 ;
        RECT 4.895000 56.540000 6.260000 57.020000 ;
        RECT 4.895000 51.100000 6.260000 51.580000 ;
        RECT 1.030000 67.420000 2.230000 67.900000 ;
        RECT 1.030000 72.860000 2.230000 73.340000 ;
        RECT 4.895000 67.420000 6.260000 67.900000 ;
        RECT 4.895000 72.860000 6.260000 73.340000 ;
        RECT 1.030000 83.740000 2.230000 84.220000 ;
        RECT 1.030000 78.300000 2.230000 78.780000 ;
        RECT 4.895000 78.300000 6.260000 78.780000 ;
        RECT 4.895000 83.740000 6.260000 84.220000 ;
        RECT 1.030000 89.180000 2.230000 89.660000 ;
        RECT 1.030000 94.620000 2.230000 95.100000 ;
        RECT 4.895000 89.180000 6.260000 89.660000 ;
        RECT 4.895000 94.620000 6.260000 95.100000 ;
        RECT 50.060000 7.580000 51.260000 8.060000 ;
        RECT 50.060000 13.020000 51.260000 13.500000 ;
        RECT 50.060000 18.460000 51.260000 18.940000 ;
        RECT 50.060000 23.900000 51.260000 24.380000 ;
        RECT 77.810000 7.580000 79.010000 8.060000 ;
        RECT 77.810000 23.900000 79.010000 24.380000 ;
        RECT 77.810000 13.020000 79.010000 13.500000 ;
        RECT 77.810000 18.460000 79.010000 18.940000 ;
        RECT 50.060000 29.340000 51.260000 29.820000 ;
        RECT 50.060000 34.780000 51.260000 35.260000 ;
        RECT 50.060000 40.220000 51.260000 40.700000 ;
        RECT 50.060000 45.660000 51.260000 46.140000 ;
        RECT 77.810000 29.340000 79.010000 29.820000 ;
        RECT 77.810000 34.780000 79.010000 35.260000 ;
        RECT 77.810000 45.660000 79.010000 46.140000 ;
        RECT 77.810000 40.220000 79.010000 40.700000 ;
        RECT 50.060000 56.540000 51.260000 57.020000 ;
        RECT 50.060000 51.100000 51.260000 51.580000 ;
        RECT 50.060000 61.980000 51.260000 62.460000 ;
        RECT 50.060000 67.420000 51.260000 67.900000 ;
        RECT 50.060000 72.860000 51.260000 73.340000 ;
        RECT 77.810000 51.100000 79.010000 51.580000 ;
        RECT 77.810000 56.540000 79.010000 57.020000 ;
        RECT 77.810000 61.980000 79.010000 62.460000 ;
        RECT 77.810000 72.860000 79.010000 73.340000 ;
        RECT 77.810000 67.420000 79.010000 67.900000 ;
        RECT 50.060000 78.300000 51.260000 78.780000 ;
        RECT 50.060000 83.740000 51.260000 84.220000 ;
        RECT 50.060000 89.180000 51.260000 89.660000 ;
        RECT 50.060000 94.620000 51.260000 95.100000 ;
        RECT 77.810000 78.300000 79.010000 78.780000 ;
        RECT 77.810000 83.740000 79.010000 84.220000 ;
        RECT 77.810000 94.620000 79.010000 95.100000 ;
        RECT 77.810000 89.180000 79.010000 89.660000 ;
        RECT 1.030000 105.500000 2.230000 105.980000 ;
        RECT 1.030000 110.940000 2.230000 111.420000 ;
        RECT 4.895000 105.500000 6.260000 105.980000 ;
        RECT 4.895000 110.940000 6.260000 111.420000 ;
        RECT 1.030000 121.820000 2.230000 122.300000 ;
        RECT 1.030000 116.380000 2.230000 116.860000 ;
        RECT 4.895000 116.380000 6.260000 116.860000 ;
        RECT 4.895000 121.820000 6.260000 122.300000 ;
        RECT 1.030000 127.260000 2.230000 127.740000 ;
        RECT 1.030000 132.700000 2.230000 133.180000 ;
        RECT 4.895000 127.260000 6.260000 127.740000 ;
        RECT 4.895000 132.700000 6.260000 133.180000 ;
        RECT 1.030000 149.020000 2.230000 149.500000 ;
        RECT 1.030000 143.580000 2.230000 144.060000 ;
        RECT 1.030000 138.140000 2.230000 138.620000 ;
        RECT 4.895000 149.020000 6.260000 149.500000 ;
        RECT 4.895000 143.580000 6.260000 144.060000 ;
        RECT 4.895000 138.140000 6.260000 138.620000 ;
        RECT 1.030000 154.460000 2.230000 154.940000 ;
        RECT 1.030000 159.900000 2.230000 160.380000 ;
        RECT 4.895000 154.460000 6.260000 154.940000 ;
        RECT 4.895000 159.900000 6.260000 160.380000 ;
        RECT 1.030000 165.340000 2.230000 165.820000 ;
        RECT 1.030000 170.780000 2.230000 171.260000 ;
        RECT 4.895000 165.340000 6.260000 165.820000 ;
        RECT 4.895000 170.780000 6.260000 171.260000 ;
        RECT 1.030000 187.100000 2.230000 187.580000 ;
        RECT 1.030000 181.660000 2.230000 182.140000 ;
        RECT 1.030000 176.220000 2.230000 176.700000 ;
        RECT 4.895000 187.100000 6.260000 187.580000 ;
        RECT 4.895000 181.660000 6.260000 182.140000 ;
        RECT 4.895000 176.220000 6.260000 176.700000 ;
        RECT 4.895000 192.540000 6.260000 193.020000 ;
        RECT 1.030000 192.540000 2.230000 193.020000 ;
        RECT 50.060000 110.940000 51.260000 111.420000 ;
        RECT 50.060000 105.500000 51.260000 105.980000 ;
        RECT 50.060000 116.380000 51.260000 116.860000 ;
        RECT 50.060000 121.820000 51.260000 122.300000 ;
        RECT 77.810000 105.500000 79.010000 105.980000 ;
        RECT 77.810000 110.940000 79.010000 111.420000 ;
        RECT 77.810000 121.820000 79.010000 122.300000 ;
        RECT 77.810000 116.380000 79.010000 116.860000 ;
        RECT 50.060000 127.260000 51.260000 127.740000 ;
        RECT 50.060000 132.700000 51.260000 133.180000 ;
        RECT 50.060000 138.140000 51.260000 138.620000 ;
        RECT 50.060000 143.580000 51.260000 144.060000 ;
        RECT 50.060000 149.020000 51.260000 149.500000 ;
        RECT 77.810000 127.260000 79.010000 127.740000 ;
        RECT 77.810000 132.700000 79.010000 133.180000 ;
        RECT 77.810000 149.020000 79.010000 149.500000 ;
        RECT 77.810000 138.140000 79.010000 138.620000 ;
        RECT 77.810000 143.580000 79.010000 144.060000 ;
        RECT 50.060000 154.460000 51.260000 154.940000 ;
        RECT 50.060000 159.900000 51.260000 160.380000 ;
        RECT 50.060000 165.340000 51.260000 165.820000 ;
        RECT 50.060000 170.780000 51.260000 171.260000 ;
        RECT 77.810000 154.460000 79.010000 154.940000 ;
        RECT 77.810000 159.900000 79.010000 160.380000 ;
        RECT 77.810000 170.780000 79.010000 171.260000 ;
        RECT 77.810000 165.340000 79.010000 165.820000 ;
        RECT 50.060000 176.220000 51.260000 176.700000 ;
        RECT 50.060000 181.660000 51.260000 182.140000 ;
        RECT 50.060000 187.100000 51.260000 187.580000 ;
        RECT 50.060000 192.540000 51.260000 193.020000 ;
        RECT 77.810000 176.220000 79.010000 176.700000 ;
        RECT 77.810000 181.660000 79.010000 182.140000 ;
        RECT 77.810000 187.100000 79.010000 187.580000 ;
        RECT 77.810000 192.540000 79.010000 193.020000 ;
      LAYER met4 ;
        RECT 50.060000 1.050000 51.260000 198.020000 ;
        RECT 5.060000 1.050000 6.260000 198.020000 ;
        RECT 77.810000 0.000000 79.010000 200.260000 ;
        RECT 1.030000 0.000000 2.230000 200.260000 ;
        RECT 4.895000 100.060000 6.260000 100.540000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 4.895000 29.340000 6.260000 29.820000 ;
        RECT 4.895000 34.780000 6.260000 35.260000 ;
        RECT 4.895000 40.220000 6.260000 40.700000 ;
        RECT 4.895000 45.660000 6.260000 46.140000 ;
        RECT 4.895000 61.980000 6.260000 62.460000 ;
        RECT 4.895000 56.540000 6.260000 57.020000 ;
        RECT 4.895000 51.100000 6.260000 51.580000 ;
        RECT 4.895000 67.420000 6.260000 67.900000 ;
        RECT 4.895000 72.860000 6.260000 73.340000 ;
        RECT 4.895000 78.300000 6.260000 78.780000 ;
        RECT 4.895000 83.740000 6.260000 84.220000 ;
        RECT 4.895000 89.180000 6.260000 89.660000 ;
        RECT 4.895000 94.620000 6.260000 95.100000 ;
        RECT 4.895000 105.500000 6.260000 105.980000 ;
        RECT 4.895000 110.940000 6.260000 111.420000 ;
        RECT 4.895000 116.380000 6.260000 116.860000 ;
        RECT 4.895000 121.820000 6.260000 122.300000 ;
        RECT 4.895000 127.260000 6.260000 127.740000 ;
        RECT 4.895000 132.700000 6.260000 133.180000 ;
        RECT 4.895000 149.020000 6.260000 149.500000 ;
        RECT 4.895000 143.580000 6.260000 144.060000 ;
        RECT 4.895000 138.140000 6.260000 138.620000 ;
        RECT 4.895000 154.460000 6.260000 154.940000 ;
        RECT 4.895000 159.900000 6.260000 160.380000 ;
        RECT 4.895000 165.340000 6.260000 165.820000 ;
        RECT 4.895000 170.780000 6.260000 171.260000 ;
        RECT 4.895000 187.100000 6.260000 187.580000 ;
        RECT 4.895000 181.660000 6.260000 182.140000 ;
        RECT 4.895000 176.220000 6.260000 176.700000 ;
        RECT 4.895000 192.540000 6.260000 193.020000 ;
    END
# end of P/G power stripe data as pin

  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 80.040000 200.260000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 80.040000 200.260000 ;
    LAYER met2 ;
      RECT 75.080000 199.420000 80.040000 200.260000 ;
      RECT 71.400000 199.420000 74.420000 200.260000 ;
      RECT 67.720000 199.420000 70.740000 200.260000 ;
      RECT 64.500000 199.420000 67.060000 200.260000 ;
      RECT 60.820000 199.420000 63.840000 200.260000 ;
      RECT 57.600000 199.420000 60.160000 200.260000 ;
      RECT 53.920000 199.420000 56.940000 200.260000 ;
      RECT 50.700000 199.420000 53.260000 200.260000 ;
      RECT 47.020000 199.420000 50.040000 200.260000 ;
      RECT 43.800000 199.420000 46.360000 200.260000 ;
      RECT 40.120000 199.420000 43.140000 200.260000 ;
      RECT 36.440000 199.420000 39.460000 200.260000 ;
      RECT 33.220000 199.420000 35.780000 200.260000 ;
      RECT 29.540000 199.420000 32.560000 200.260000 ;
      RECT 26.320000 199.420000 28.880000 200.260000 ;
      RECT 22.640000 199.420000 25.660000 200.260000 ;
      RECT 19.420000 199.420000 21.980000 200.260000 ;
      RECT 15.740000 199.420000 18.760000 200.260000 ;
      RECT 12.520000 199.420000 15.080000 200.260000 ;
      RECT 8.840000 199.420000 11.860000 200.260000 ;
      RECT 5.620000 199.420000 8.180000 200.260000 ;
      RECT 0.000000 199.420000 4.960000 200.260000 ;
      RECT 0.000000 0.840000 80.040000 199.420000 ;
      RECT 75.080000 0.000000 80.040000 0.840000 ;
      RECT 71.400000 0.000000 74.420000 0.840000 ;
      RECT 67.720000 0.000000 70.740000 0.840000 ;
      RECT 64.500000 0.000000 67.060000 0.840000 ;
      RECT 60.820000 0.000000 63.840000 0.840000 ;
      RECT 57.600000 0.000000 60.160000 0.840000 ;
      RECT 53.920000 0.000000 56.940000 0.840000 ;
      RECT 50.700000 0.000000 53.260000 0.840000 ;
      RECT 47.020000 0.000000 50.040000 0.840000 ;
      RECT 43.800000 0.000000 46.360000 0.840000 ;
      RECT 40.120000 0.000000 43.140000 0.840000 ;
      RECT 36.440000 0.000000 39.460000 0.840000 ;
      RECT 33.220000 0.000000 35.780000 0.840000 ;
      RECT 29.540000 0.000000 32.560000 0.840000 ;
      RECT 26.320000 0.000000 28.880000 0.840000 ;
      RECT 22.640000 0.000000 25.660000 0.840000 ;
      RECT 19.420000 0.000000 21.980000 0.840000 ;
      RECT 15.740000 0.000000 18.760000 0.840000 ;
      RECT 12.520000 0.000000 15.080000 0.840000 ;
      RECT 8.840000 0.000000 11.860000 0.840000 ;
      RECT 5.620000 0.000000 8.180000 0.840000 ;
      RECT 0.000000 0.000000 4.960000 0.840000 ;
    LAYER met3 ;
      RECT 0.000000 198.320000 80.040000 200.260000 ;
      RECT 1.000000 193.880000 79.040000 194.720000 ;
      RECT 0.000000 193.320000 80.040000 193.880000 ;
      RECT 79.310000 193.030000 80.040000 193.320000 ;
      RECT 51.560000 192.240000 77.510000 193.320000 ;
      RECT 6.560000 192.240000 49.760000 193.320000 ;
      RECT 2.530000 192.240000 4.595000 193.320000 ;
      RECT 0.000000 192.240000 0.730000 193.320000 ;
      RECT 0.000000 192.050000 79.040000 192.240000 ;
      RECT 0.000000 191.810000 80.040000 192.050000 ;
      RECT 0.000000 190.830000 79.040000 191.810000 ;
      RECT 0.000000 190.600000 80.040000 190.830000 ;
      RECT 0.000000 190.590000 2.530000 190.600000 ;
      RECT 77.510000 189.980000 80.040000 190.600000 ;
      RECT 1.000000 189.610000 2.530000 190.590000 ;
      RECT 77.510000 189.520000 79.040000 189.980000 ;
      RECT 53.560000 189.520000 75.710000 190.600000 ;
      RECT 8.560000 189.520000 51.760000 190.600000 ;
      RECT 4.330000 189.520000 6.760000 190.600000 ;
      RECT 0.000000 189.520000 2.530000 189.610000 ;
      RECT 0.000000 189.000000 79.040000 189.520000 ;
      RECT 0.000000 188.760000 80.040000 189.000000 ;
      RECT 0.000000 187.880000 79.040000 188.760000 ;
      RECT 79.310000 186.930000 80.040000 187.780000 ;
      RECT 51.560000 186.800000 77.510000 187.880000 ;
      RECT 6.560000 186.800000 49.760000 187.880000 ;
      RECT 2.530000 186.800000 4.595000 187.880000 ;
      RECT 0.000000 186.800000 0.730000 187.880000 ;
      RECT 0.000000 186.320000 79.040000 186.800000 ;
      RECT 1.000000 185.950000 79.040000 186.320000 ;
      RECT 1.000000 185.710000 80.040000 185.950000 ;
      RECT 1.000000 185.340000 79.040000 185.710000 ;
      RECT 0.000000 185.160000 79.040000 185.340000 ;
      RECT 77.510000 184.730000 79.040000 185.160000 ;
      RECT 77.510000 184.080000 80.040000 184.730000 ;
      RECT 53.560000 184.080000 75.710000 185.160000 ;
      RECT 8.560000 184.080000 51.760000 185.160000 ;
      RECT 4.330000 184.080000 6.760000 185.160000 ;
      RECT 0.000000 184.080000 2.530000 185.160000 ;
      RECT 0.000000 183.880000 80.040000 184.080000 ;
      RECT 0.000000 182.900000 79.040000 183.880000 ;
      RECT 0.000000 182.660000 80.040000 182.900000 ;
      RECT 0.000000 182.440000 79.040000 182.660000 ;
      RECT 0.000000 182.050000 0.730000 182.440000 ;
      RECT 79.310000 181.440000 80.040000 181.680000 ;
      RECT 51.560000 181.360000 77.510000 182.440000 ;
      RECT 6.560000 181.360000 49.760000 182.440000 ;
      RECT 2.530000 181.360000 4.595000 182.440000 ;
      RECT 1.000000 181.070000 79.040000 181.360000 ;
      RECT 0.000000 180.460000 79.040000 181.070000 ;
      RECT 0.000000 179.720000 80.040000 180.460000 ;
      RECT 77.510000 179.610000 80.040000 179.720000 ;
      RECT 77.510000 178.640000 79.040000 179.610000 ;
      RECT 53.560000 178.640000 75.710000 179.720000 ;
      RECT 8.560000 178.640000 51.760000 179.720000 ;
      RECT 4.330000 178.640000 6.760000 179.720000 ;
      RECT 0.000000 178.640000 2.530000 179.720000 ;
      RECT 0.000000 178.630000 79.040000 178.640000 ;
      RECT 0.000000 178.390000 80.040000 178.630000 ;
      RECT 0.000000 177.780000 79.040000 178.390000 ;
      RECT 1.000000 177.410000 79.040000 177.780000 ;
      RECT 1.000000 177.000000 80.040000 177.410000 ;
      RECT 79.310000 176.560000 80.040000 177.000000 ;
      RECT 51.560000 175.920000 77.510000 177.000000 ;
      RECT 6.560000 175.920000 49.760000 177.000000 ;
      RECT 2.530000 175.920000 4.595000 177.000000 ;
      RECT 0.000000 175.920000 0.730000 176.800000 ;
      RECT 0.000000 175.580000 79.040000 175.920000 ;
      RECT 0.000000 175.340000 80.040000 175.580000 ;
      RECT 0.000000 174.360000 79.040000 175.340000 ;
      RECT 0.000000 174.280000 80.040000 174.360000 ;
      RECT 77.510000 173.510000 80.040000 174.280000 ;
      RECT 0.000000 173.510000 2.530000 174.280000 ;
      RECT 77.510000 173.200000 79.040000 173.510000 ;
      RECT 53.560000 173.200000 75.710000 174.280000 ;
      RECT 8.560000 173.200000 51.760000 174.280000 ;
      RECT 4.330000 173.200000 6.760000 174.280000 ;
      RECT 1.000000 173.200000 2.530000 173.510000 ;
      RECT 1.000000 172.530000 79.040000 173.200000 ;
      RECT 0.000000 172.290000 80.040000 172.530000 ;
      RECT 0.000000 171.560000 79.040000 172.290000 ;
      RECT 79.310000 170.480000 80.040000 171.310000 ;
      RECT 51.560000 170.480000 77.510000 171.560000 ;
      RECT 6.560000 170.480000 49.760000 171.560000 ;
      RECT 2.530000 170.480000 4.595000 171.560000 ;
      RECT 0.000000 170.480000 0.730000 171.560000 ;
      RECT 0.000000 170.460000 80.040000 170.480000 ;
      RECT 0.000000 169.480000 79.040000 170.460000 ;
      RECT 0.000000 169.240000 80.040000 169.480000 ;
      RECT 1.000000 168.840000 79.040000 169.240000 ;
      RECT 77.510000 168.260000 79.040000 168.840000 ;
      RECT 1.000000 168.260000 2.530000 168.840000 ;
      RECT 77.510000 168.020000 80.040000 168.260000 ;
      RECT 77.510000 167.760000 79.040000 168.020000 ;
      RECT 53.560000 167.760000 75.710000 168.840000 ;
      RECT 8.560000 167.760000 51.760000 168.840000 ;
      RECT 4.330000 167.760000 6.760000 168.840000 ;
      RECT 0.000000 167.760000 2.530000 168.260000 ;
      RECT 0.000000 167.040000 79.040000 167.760000 ;
      RECT 0.000000 166.190000 80.040000 167.040000 ;
      RECT 0.000000 166.120000 79.040000 166.190000 ;
      RECT 79.310000 165.040000 80.040000 165.210000 ;
      RECT 51.560000 165.040000 77.510000 166.120000 ;
      RECT 6.560000 165.040000 49.760000 166.120000 ;
      RECT 2.530000 165.040000 4.595000 166.120000 ;
      RECT 0.000000 165.040000 0.730000 166.120000 ;
      RECT 0.000000 164.970000 80.040000 165.040000 ;
      RECT 1.000000 163.990000 79.040000 164.970000 ;
      RECT 0.000000 163.400000 80.040000 163.990000 ;
      RECT 77.510000 163.140000 80.040000 163.400000 ;
      RECT 77.510000 162.320000 79.040000 163.140000 ;
      RECT 53.560000 162.320000 75.710000 163.400000 ;
      RECT 8.560000 162.320000 51.760000 163.400000 ;
      RECT 4.330000 162.320000 6.760000 163.400000 ;
      RECT 0.000000 162.320000 2.530000 163.400000 ;
      RECT 0.000000 162.160000 79.040000 162.320000 ;
      RECT 0.000000 161.920000 80.040000 162.160000 ;
      RECT 0.000000 160.940000 79.040000 161.920000 ;
      RECT 0.000000 160.700000 80.040000 160.940000 ;
      RECT 1.000000 160.680000 80.040000 160.700000 ;
      RECT 79.310000 160.090000 80.040000 160.680000 ;
      RECT 51.560000 159.600000 77.510000 160.680000 ;
      RECT 6.560000 159.600000 49.760000 160.680000 ;
      RECT 2.530000 159.600000 4.595000 160.680000 ;
      RECT 0.000000 159.600000 0.730000 159.720000 ;
      RECT 0.000000 159.110000 79.040000 159.600000 ;
      RECT 0.000000 158.870000 80.040000 159.110000 ;
      RECT 0.000000 157.960000 79.040000 158.870000 ;
      RECT 77.510000 157.890000 79.040000 157.960000 ;
      RECT 77.510000 157.040000 80.040000 157.890000 ;
      RECT 77.510000 156.880000 79.040000 157.040000 ;
      RECT 53.560000 156.880000 75.710000 157.960000 ;
      RECT 8.560000 156.880000 51.760000 157.960000 ;
      RECT 4.330000 156.880000 6.760000 157.960000 ;
      RECT 0.000000 156.880000 2.530000 157.960000 ;
      RECT 0.000000 156.430000 79.040000 156.880000 ;
      RECT 1.000000 156.060000 79.040000 156.430000 ;
      RECT 1.000000 155.820000 80.040000 156.060000 ;
      RECT 1.000000 155.450000 79.040000 155.820000 ;
      RECT 0.000000 155.240000 79.040000 155.450000 ;
      RECT 79.310000 154.600000 80.040000 154.840000 ;
      RECT 51.560000 154.160000 77.510000 155.240000 ;
      RECT 6.560000 154.160000 49.760000 155.240000 ;
      RECT 2.530000 154.160000 4.595000 155.240000 ;
      RECT 0.000000 154.160000 0.730000 155.240000 ;
      RECT 0.000000 153.620000 79.040000 154.160000 ;
      RECT 0.000000 152.770000 80.040000 153.620000 ;
      RECT 1.000000 152.520000 79.040000 152.770000 ;
      RECT 77.510000 151.790000 79.040000 152.520000 ;
      RECT 1.000000 151.790000 2.530000 152.520000 ;
      RECT 77.510000 151.550000 80.040000 151.790000 ;
      RECT 77.510000 151.440000 79.040000 151.550000 ;
      RECT 53.560000 151.440000 75.710000 152.520000 ;
      RECT 8.560000 151.440000 51.760000 152.520000 ;
      RECT 4.330000 151.440000 6.760000 152.520000 ;
      RECT 0.000000 151.440000 2.530000 151.790000 ;
      RECT 0.000000 150.570000 79.040000 151.440000 ;
      RECT 0.000000 149.800000 80.040000 150.570000 ;
      RECT 79.310000 149.720000 80.040000 149.800000 ;
      RECT 79.310000 148.720000 80.040000 148.740000 ;
      RECT 51.560000 148.720000 77.510000 149.800000 ;
      RECT 6.560000 148.720000 49.760000 149.800000 ;
      RECT 2.530000 148.720000 4.595000 149.800000 ;
      RECT 0.000000 148.720000 0.730000 149.800000 ;
      RECT 0.000000 148.500000 80.040000 148.720000 ;
      RECT 1.000000 147.520000 79.040000 148.500000 ;
      RECT 0.000000 147.080000 80.040000 147.520000 ;
      RECT 77.510000 146.670000 80.040000 147.080000 ;
      RECT 77.510000 146.000000 79.040000 146.670000 ;
      RECT 53.560000 146.000000 75.710000 147.080000 ;
      RECT 8.560000 146.000000 51.760000 147.080000 ;
      RECT 4.330000 146.000000 6.760000 147.080000 ;
      RECT 0.000000 146.000000 2.530000 147.080000 ;
      RECT 0.000000 145.690000 79.040000 146.000000 ;
      RECT 0.000000 145.450000 80.040000 145.690000 ;
      RECT 0.000000 144.470000 79.040000 145.450000 ;
      RECT 0.000000 144.360000 80.040000 144.470000 ;
      RECT 79.310000 144.230000 80.040000 144.360000 ;
      RECT 0.000000 144.230000 0.730000 144.360000 ;
      RECT 51.560000 143.280000 77.510000 144.360000 ;
      RECT 6.560000 143.280000 49.760000 144.360000 ;
      RECT 2.530000 143.280000 4.595000 144.360000 ;
      RECT 1.000000 143.250000 79.040000 143.280000 ;
      RECT 0.000000 142.400000 80.040000 143.250000 ;
      RECT 0.000000 141.640000 79.040000 142.400000 ;
      RECT 77.510000 141.420000 79.040000 141.640000 ;
      RECT 77.510000 141.180000 80.040000 141.420000 ;
      RECT 77.510000 140.560000 79.040000 141.180000 ;
      RECT 53.560000 140.560000 75.710000 141.640000 ;
      RECT 8.560000 140.560000 51.760000 141.640000 ;
      RECT 4.330000 140.560000 6.760000 141.640000 ;
      RECT 0.000000 140.560000 2.530000 141.640000 ;
      RECT 0.000000 140.200000 79.040000 140.560000 ;
      RECT 0.000000 139.960000 80.040000 140.200000 ;
      RECT 1.000000 139.350000 80.040000 139.960000 ;
      RECT 1.000000 138.980000 79.040000 139.350000 ;
      RECT 0.000000 138.920000 79.040000 138.980000 ;
      RECT 79.310000 138.130000 80.040000 138.370000 ;
      RECT 51.560000 137.840000 77.510000 138.920000 ;
      RECT 6.560000 137.840000 49.760000 138.920000 ;
      RECT 2.530000 137.840000 4.595000 138.920000 ;
      RECT 0.000000 137.840000 0.730000 138.920000 ;
      RECT 0.000000 137.150000 79.040000 137.840000 ;
      RECT 0.000000 136.300000 80.040000 137.150000 ;
      RECT 0.000000 136.200000 79.040000 136.300000 ;
      RECT 0.000000 135.690000 2.530000 136.200000 ;
      RECT 77.510000 135.320000 79.040000 136.200000 ;
      RECT 77.510000 135.120000 80.040000 135.320000 ;
      RECT 53.560000 135.120000 75.710000 136.200000 ;
      RECT 8.560000 135.120000 51.760000 136.200000 ;
      RECT 4.330000 135.120000 6.760000 136.200000 ;
      RECT 1.000000 135.120000 2.530000 135.690000 ;
      RECT 1.000000 135.080000 80.040000 135.120000 ;
      RECT 1.000000 134.710000 79.040000 135.080000 ;
      RECT 0.000000 134.100000 79.040000 134.710000 ;
      RECT 0.000000 133.480000 80.040000 134.100000 ;
      RECT 79.310000 133.250000 80.040000 133.480000 ;
      RECT 51.560000 132.400000 77.510000 133.480000 ;
      RECT 6.560000 132.400000 49.760000 133.480000 ;
      RECT 2.530000 132.400000 4.595000 133.480000 ;
      RECT 0.000000 132.400000 0.730000 133.480000 ;
      RECT 0.000000 132.270000 79.040000 132.400000 ;
      RECT 0.000000 132.030000 80.040000 132.270000 ;
      RECT 0.000000 131.420000 79.040000 132.030000 ;
      RECT 1.000000 131.050000 79.040000 131.420000 ;
      RECT 1.000000 130.810000 80.040000 131.050000 ;
      RECT 1.000000 130.760000 79.040000 130.810000 ;
      RECT 1.000000 130.440000 2.530000 130.760000 ;
      RECT 77.510000 129.830000 79.040000 130.760000 ;
      RECT 77.510000 129.680000 80.040000 129.830000 ;
      RECT 53.560000 129.680000 75.710000 130.760000 ;
      RECT 8.560000 129.680000 51.760000 130.760000 ;
      RECT 4.330000 129.680000 6.760000 130.760000 ;
      RECT 0.000000 129.680000 2.530000 130.440000 ;
      RECT 0.000000 128.980000 80.040000 129.680000 ;
      RECT 0.000000 128.040000 79.040000 128.980000 ;
      RECT 79.310000 127.760000 80.040000 128.000000 ;
      RECT 0.000000 127.150000 0.730000 128.040000 ;
      RECT 51.560000 126.960000 77.510000 128.040000 ;
      RECT 6.560000 126.960000 49.760000 128.040000 ;
      RECT 2.530000 126.960000 4.595000 128.040000 ;
      RECT 1.000000 126.780000 79.040000 126.960000 ;
      RECT 1.000000 126.170000 80.040000 126.780000 ;
      RECT 0.000000 125.930000 80.040000 126.170000 ;
      RECT 0.000000 125.320000 79.040000 125.930000 ;
      RECT 77.510000 124.950000 79.040000 125.320000 ;
      RECT 77.510000 124.710000 80.040000 124.950000 ;
      RECT 77.510000 124.240000 79.040000 124.710000 ;
      RECT 53.560000 124.240000 75.710000 125.320000 ;
      RECT 8.560000 124.240000 51.760000 125.320000 ;
      RECT 4.330000 124.240000 6.760000 125.320000 ;
      RECT 0.000000 124.240000 2.530000 125.320000 ;
      RECT 0.000000 123.730000 79.040000 124.240000 ;
      RECT 0.000000 122.880000 80.040000 123.730000 ;
      RECT 1.000000 122.600000 79.040000 122.880000 ;
      RECT 79.310000 121.660000 80.040000 121.900000 ;
      RECT 51.560000 121.520000 77.510000 122.600000 ;
      RECT 6.560000 121.520000 49.760000 122.600000 ;
      RECT 2.530000 121.520000 4.595000 122.600000 ;
      RECT 0.000000 121.520000 0.730000 121.900000 ;
      RECT 0.000000 120.680000 79.040000 121.520000 ;
      RECT 0.000000 119.880000 80.040000 120.680000 ;
      RECT 77.510000 119.830000 80.040000 119.880000 ;
      RECT 77.510000 118.850000 79.040000 119.830000 ;
      RECT 77.510000 118.800000 80.040000 118.850000 ;
      RECT 53.560000 118.800000 75.710000 119.880000 ;
      RECT 8.560000 118.800000 51.760000 119.880000 ;
      RECT 4.330000 118.800000 6.760000 119.880000 ;
      RECT 0.000000 118.800000 2.530000 119.880000 ;
      RECT 0.000000 118.610000 80.040000 118.800000 ;
      RECT 1.000000 117.630000 79.040000 118.610000 ;
      RECT 0.000000 117.390000 80.040000 117.630000 ;
      RECT 0.000000 117.160000 79.040000 117.390000 ;
      RECT 79.310000 116.080000 80.040000 116.410000 ;
      RECT 51.560000 116.080000 77.510000 117.160000 ;
      RECT 6.560000 116.080000 49.760000 117.160000 ;
      RECT 2.530000 116.080000 4.595000 117.160000 ;
      RECT 0.000000 116.080000 0.730000 117.160000 ;
      RECT 0.000000 115.560000 80.040000 116.080000 ;
      RECT 0.000000 114.950000 79.040000 115.560000 ;
      RECT 1.000000 114.580000 79.040000 114.950000 ;
      RECT 1.000000 114.440000 80.040000 114.580000 ;
      RECT 77.510000 114.340000 80.040000 114.440000 ;
      RECT 1.000000 113.970000 2.530000 114.440000 ;
      RECT 77.510000 113.360000 79.040000 114.340000 ;
      RECT 53.560000 113.360000 75.710000 114.440000 ;
      RECT 8.560000 113.360000 51.760000 114.440000 ;
      RECT 4.330000 113.360000 6.760000 114.440000 ;
      RECT 0.000000 113.360000 2.530000 113.970000 ;
      RECT 0.000000 112.510000 80.040000 113.360000 ;
      RECT 0.000000 111.720000 79.040000 112.510000 ;
      RECT 79.310000 111.290000 80.040000 111.530000 ;
      RECT 0.000000 110.680000 0.730000 111.720000 ;
      RECT 51.560000 110.640000 77.510000 111.720000 ;
      RECT 6.560000 110.640000 49.760000 111.720000 ;
      RECT 2.530000 110.640000 4.595000 111.720000 ;
      RECT 1.000000 110.310000 79.040000 110.640000 ;
      RECT 1.000000 109.700000 80.040000 110.310000 ;
      RECT 0.000000 109.460000 80.040000 109.700000 ;
      RECT 0.000000 109.000000 79.040000 109.460000 ;
      RECT 77.510000 108.480000 79.040000 109.000000 ;
      RECT 77.510000 108.240000 80.040000 108.480000 ;
      RECT 77.510000 107.920000 79.040000 108.240000 ;
      RECT 53.560000 107.920000 75.710000 109.000000 ;
      RECT 8.560000 107.920000 51.760000 109.000000 ;
      RECT 4.330000 107.920000 6.760000 109.000000 ;
      RECT 0.000000 107.920000 2.530000 109.000000 ;
      RECT 0.000000 107.260000 79.040000 107.920000 ;
      RECT 0.000000 106.410000 80.040000 107.260000 ;
      RECT 1.000000 106.280000 79.040000 106.410000 ;
      RECT 79.310000 105.200000 80.040000 105.430000 ;
      RECT 51.560000 105.200000 77.510000 106.280000 ;
      RECT 6.560000 105.200000 49.760000 106.280000 ;
      RECT 2.530000 105.200000 4.595000 106.280000 ;
      RECT 0.000000 105.200000 0.730000 105.430000 ;
      RECT 0.000000 105.190000 80.040000 105.200000 ;
      RECT 0.000000 104.210000 79.040000 105.190000 ;
      RECT 0.000000 103.970000 80.040000 104.210000 ;
      RECT 0.000000 103.560000 79.040000 103.970000 ;
      RECT 77.510000 102.990000 79.040000 103.560000 ;
      RECT 77.510000 102.480000 80.040000 102.990000 ;
      RECT 53.560000 102.480000 75.710000 103.560000 ;
      RECT 8.560000 102.480000 51.760000 103.560000 ;
      RECT 4.330000 102.480000 6.760000 103.560000 ;
      RECT 0.000000 102.480000 2.530000 103.560000 ;
      RECT 0.000000 102.140000 80.040000 102.480000 ;
      RECT 1.000000 101.160000 79.040000 102.140000 ;
      RECT 0.000000 100.920000 80.040000 101.160000 ;
      RECT 0.000000 100.840000 79.040000 100.920000 ;
      RECT 79.310000 99.760000 80.040000 99.940000 ;
      RECT 51.560000 99.760000 77.510000 100.840000 ;
      RECT 6.560000 99.760000 49.760000 100.840000 ;
      RECT 2.530000 99.760000 4.595000 100.840000 ;
      RECT 0.000000 99.760000 0.730000 100.840000 ;
      RECT 0.000000 99.090000 80.040000 99.760000 ;
      RECT 0.000000 98.120000 79.040000 99.090000 ;
      RECT 77.510000 98.110000 79.040000 98.120000 ;
      RECT 77.510000 97.870000 80.040000 98.110000 ;
      RECT 0.000000 97.870000 2.530000 98.120000 ;
      RECT 77.510000 97.040000 79.040000 97.870000 ;
      RECT 53.560000 97.040000 75.710000 98.120000 ;
      RECT 8.560000 97.040000 51.760000 98.120000 ;
      RECT 4.330000 97.040000 6.760000 98.120000 ;
      RECT 1.000000 97.040000 2.530000 97.870000 ;
      RECT 1.000000 96.890000 79.040000 97.040000 ;
      RECT 0.000000 96.040000 80.040000 96.890000 ;
      RECT 0.000000 95.400000 79.040000 96.040000 ;
      RECT 79.310000 94.820000 80.040000 95.060000 ;
      RECT 51.560000 94.320000 77.510000 95.400000 ;
      RECT 6.560000 94.320000 49.760000 95.400000 ;
      RECT 2.530000 94.320000 4.595000 95.400000 ;
      RECT 0.000000 94.320000 0.730000 95.400000 ;
      RECT 0.000000 93.840000 79.040000 94.320000 ;
      RECT 0.000000 93.600000 80.040000 93.840000 ;
      RECT 1.000000 92.680000 79.040000 93.600000 ;
      RECT 77.510000 92.620000 79.040000 92.680000 ;
      RECT 1.000000 92.620000 2.530000 92.680000 ;
      RECT 77.510000 91.770000 80.040000 92.620000 ;
      RECT 77.510000 91.600000 79.040000 91.770000 ;
      RECT 53.560000 91.600000 75.710000 92.680000 ;
      RECT 8.560000 91.600000 51.760000 92.680000 ;
      RECT 4.330000 91.600000 6.760000 92.680000 ;
      RECT 0.000000 91.600000 2.530000 92.620000 ;
      RECT 0.000000 90.790000 79.040000 91.600000 ;
      RECT 0.000000 90.550000 80.040000 90.790000 ;
      RECT 0.000000 89.960000 79.040000 90.550000 ;
      RECT 0.000000 89.330000 0.730000 89.960000 ;
      RECT 79.310000 88.880000 80.040000 89.570000 ;
      RECT 51.560000 88.880000 77.510000 89.960000 ;
      RECT 6.560000 88.880000 49.760000 89.960000 ;
      RECT 2.530000 88.880000 4.595000 89.960000 ;
      RECT 1.000000 88.720000 80.040000 88.880000 ;
      RECT 1.000000 88.350000 79.040000 88.720000 ;
      RECT 0.000000 87.740000 79.040000 88.350000 ;
      RECT 0.000000 87.500000 80.040000 87.740000 ;
      RECT 0.000000 87.240000 79.040000 87.500000 ;
      RECT 77.510000 86.520000 79.040000 87.240000 ;
      RECT 77.510000 86.160000 80.040000 86.520000 ;
      RECT 53.560000 86.160000 75.710000 87.240000 ;
      RECT 8.560000 86.160000 51.760000 87.240000 ;
      RECT 4.330000 86.160000 6.760000 87.240000 ;
      RECT 0.000000 86.160000 2.530000 87.240000 ;
      RECT 0.000000 85.670000 80.040000 86.160000 ;
      RECT 0.000000 85.060000 79.040000 85.670000 ;
      RECT 1.000000 84.690000 79.040000 85.060000 ;
      RECT 1.000000 84.520000 80.040000 84.690000 ;
      RECT 79.310000 84.450000 80.040000 84.520000 ;
      RECT 79.310000 83.440000 80.040000 83.470000 ;
      RECT 51.560000 83.440000 77.510000 84.520000 ;
      RECT 6.560000 83.440000 49.760000 84.520000 ;
      RECT 2.530000 83.440000 4.595000 84.520000 ;
      RECT 0.000000 83.440000 0.730000 84.080000 ;
      RECT 0.000000 82.620000 80.040000 83.440000 ;
      RECT 0.000000 81.800000 79.040000 82.620000 ;
      RECT 77.510000 81.640000 79.040000 81.800000 ;
      RECT 77.510000 81.400000 80.040000 81.640000 ;
      RECT 0.000000 80.790000 2.530000 81.800000 ;
      RECT 77.510000 80.720000 79.040000 81.400000 ;
      RECT 53.560000 80.720000 75.710000 81.800000 ;
      RECT 8.560000 80.720000 51.760000 81.800000 ;
      RECT 4.330000 80.720000 6.760000 81.800000 ;
      RECT 1.000000 80.720000 2.530000 80.790000 ;
      RECT 1.000000 80.420000 79.040000 80.720000 ;
      RECT 1.000000 80.180000 80.040000 80.420000 ;
      RECT 1.000000 79.810000 79.040000 80.180000 ;
      RECT 0.000000 79.200000 79.040000 79.810000 ;
      RECT 0.000000 79.080000 80.040000 79.200000 ;
      RECT 79.310000 78.350000 80.040000 79.080000 ;
      RECT 51.560000 78.000000 77.510000 79.080000 ;
      RECT 6.560000 78.000000 49.760000 79.080000 ;
      RECT 2.530000 78.000000 4.595000 79.080000 ;
      RECT 0.000000 78.000000 0.730000 79.080000 ;
      RECT 0.000000 77.370000 79.040000 78.000000 ;
      RECT 0.000000 77.130000 80.040000 77.370000 ;
      RECT 1.000000 76.360000 79.040000 77.130000 ;
      RECT 77.510000 76.150000 79.040000 76.360000 ;
      RECT 1.000000 76.150000 2.530000 76.360000 ;
      RECT 77.510000 75.300000 80.040000 76.150000 ;
      RECT 77.510000 75.280000 79.040000 75.300000 ;
      RECT 53.560000 75.280000 75.710000 76.360000 ;
      RECT 8.560000 75.280000 51.760000 76.360000 ;
      RECT 4.330000 75.280000 6.760000 76.360000 ;
      RECT 0.000000 75.280000 2.530000 76.150000 ;
      RECT 0.000000 74.320000 79.040000 75.280000 ;
      RECT 0.000000 74.080000 80.040000 74.320000 ;
      RECT 0.000000 73.640000 79.040000 74.080000 ;
      RECT 0.000000 72.860000 0.730000 73.640000 ;
      RECT 79.310000 72.560000 80.040000 73.100000 ;
      RECT 51.560000 72.560000 77.510000 73.640000 ;
      RECT 6.560000 72.560000 49.760000 73.640000 ;
      RECT 2.530000 72.560000 4.595000 73.640000 ;
      RECT 1.000000 72.250000 80.040000 72.560000 ;
      RECT 1.000000 71.880000 79.040000 72.250000 ;
      RECT 0.000000 71.270000 79.040000 71.880000 ;
      RECT 0.000000 71.030000 80.040000 71.270000 ;
      RECT 0.000000 70.920000 79.040000 71.030000 ;
      RECT 77.510000 70.050000 79.040000 70.920000 ;
      RECT 77.510000 69.840000 80.040000 70.050000 ;
      RECT 53.560000 69.840000 75.710000 70.920000 ;
      RECT 8.560000 69.840000 51.760000 70.920000 ;
      RECT 4.330000 69.840000 6.760000 70.920000 ;
      RECT 0.000000 69.840000 2.530000 70.920000 ;
      RECT 0.000000 69.200000 80.040000 69.840000 ;
      RECT 0.000000 68.590000 79.040000 69.200000 ;
      RECT 1.000000 68.220000 79.040000 68.590000 ;
      RECT 1.000000 68.200000 80.040000 68.220000 ;
      RECT 79.310000 67.980000 80.040000 68.200000 ;
      RECT 51.560000 67.120000 77.510000 68.200000 ;
      RECT 6.560000 67.120000 49.760000 68.200000 ;
      RECT 2.530000 67.120000 4.595000 68.200000 ;
      RECT 0.000000 67.120000 0.730000 67.610000 ;
      RECT 0.000000 67.000000 79.040000 67.120000 ;
      RECT 0.000000 66.760000 80.040000 67.000000 ;
      RECT 0.000000 65.780000 79.040000 66.760000 ;
      RECT 0.000000 65.480000 80.040000 65.780000 ;
      RECT 77.510000 64.930000 80.040000 65.480000 ;
      RECT 77.510000 64.400000 79.040000 64.930000 ;
      RECT 53.560000 64.400000 75.710000 65.480000 ;
      RECT 8.560000 64.400000 51.760000 65.480000 ;
      RECT 4.330000 64.400000 6.760000 65.480000 ;
      RECT 0.000000 64.400000 2.530000 65.480000 ;
      RECT 0.000000 64.320000 79.040000 64.400000 ;
      RECT 1.000000 63.950000 79.040000 64.320000 ;
      RECT 1.000000 63.710000 80.040000 63.950000 ;
      RECT 1.000000 63.340000 79.040000 63.710000 ;
      RECT 0.000000 62.760000 79.040000 63.340000 ;
      RECT 79.310000 61.880000 80.040000 62.730000 ;
      RECT 51.560000 61.680000 77.510000 62.760000 ;
      RECT 6.560000 61.680000 49.760000 62.760000 ;
      RECT 2.530000 61.680000 4.595000 62.760000 ;
      RECT 0.000000 61.680000 0.730000 62.760000 ;
      RECT 0.000000 60.900000 79.040000 61.680000 ;
      RECT 0.000000 60.660000 80.040000 60.900000 ;
      RECT 0.000000 60.050000 79.040000 60.660000 ;
      RECT 1.000000 60.040000 79.040000 60.050000 ;
      RECT 77.510000 59.680000 79.040000 60.040000 ;
      RECT 1.000000 59.070000 2.530000 60.040000 ;
      RECT 77.510000 58.960000 80.040000 59.680000 ;
      RECT 53.560000 58.960000 75.710000 60.040000 ;
      RECT 8.560000 58.960000 51.760000 60.040000 ;
      RECT 4.330000 58.960000 6.760000 60.040000 ;
      RECT 0.000000 58.960000 2.530000 59.070000 ;
      RECT 0.000000 58.830000 80.040000 58.960000 ;
      RECT 0.000000 57.850000 79.040000 58.830000 ;
      RECT 0.000000 57.610000 80.040000 57.850000 ;
      RECT 0.000000 57.320000 79.040000 57.610000 ;
      RECT 79.310000 56.240000 80.040000 56.630000 ;
      RECT 51.560000 56.240000 77.510000 57.320000 ;
      RECT 6.560000 56.240000 49.760000 57.320000 ;
      RECT 2.530000 56.240000 4.595000 57.320000 ;
      RECT 0.000000 56.240000 0.730000 57.320000 ;
      RECT 0.000000 55.780000 80.040000 56.240000 ;
      RECT 1.000000 54.800000 79.040000 55.780000 ;
      RECT 0.000000 54.600000 80.040000 54.800000 ;
      RECT 77.510000 54.560000 80.040000 54.600000 ;
      RECT 77.510000 53.580000 79.040000 54.560000 ;
      RECT 77.510000 53.520000 80.040000 53.580000 ;
      RECT 53.560000 53.520000 75.710000 54.600000 ;
      RECT 8.560000 53.520000 51.760000 54.600000 ;
      RECT 4.330000 53.520000 6.760000 54.600000 ;
      RECT 0.000000 53.520000 2.530000 54.600000 ;
      RECT 0.000000 53.340000 80.040000 53.520000 ;
      RECT 0.000000 52.360000 79.040000 53.340000 ;
      RECT 0.000000 51.880000 80.040000 52.360000 ;
      RECT 79.310000 51.510000 80.040000 51.880000 ;
      RECT 0.000000 51.510000 0.730000 51.880000 ;
      RECT 51.560000 50.800000 77.510000 51.880000 ;
      RECT 6.560000 50.800000 49.760000 51.880000 ;
      RECT 2.530000 50.800000 4.595000 51.880000 ;
      RECT 1.000000 50.530000 79.040000 50.800000 ;
      RECT 0.000000 50.290000 80.040000 50.530000 ;
      RECT 0.000000 49.310000 79.040000 50.290000 ;
      RECT 0.000000 49.160000 80.040000 49.310000 ;
      RECT 77.510000 48.460000 80.040000 49.160000 ;
      RECT 77.510000 48.080000 79.040000 48.460000 ;
      RECT 53.560000 48.080000 75.710000 49.160000 ;
      RECT 8.560000 48.080000 51.760000 49.160000 ;
      RECT 4.330000 48.080000 6.760000 49.160000 ;
      RECT 0.000000 48.080000 2.530000 49.160000 ;
      RECT 0.000000 47.480000 79.040000 48.080000 ;
      RECT 0.000000 47.240000 80.040000 47.480000 ;
      RECT 1.000000 46.440000 79.040000 47.240000 ;
      RECT 79.310000 45.410000 80.040000 46.260000 ;
      RECT 51.560000 45.360000 77.510000 46.440000 ;
      RECT 6.560000 45.360000 49.760000 46.440000 ;
      RECT 2.530000 45.360000 4.595000 46.440000 ;
      RECT 0.000000 45.360000 0.730000 46.260000 ;
      RECT 0.000000 44.430000 79.040000 45.360000 ;
      RECT 0.000000 44.190000 80.040000 44.430000 ;
      RECT 0.000000 43.720000 79.040000 44.190000 ;
      RECT 77.510000 43.210000 79.040000 43.720000 ;
      RECT 77.510000 42.970000 80.040000 43.210000 ;
      RECT 0.000000 42.970000 2.530000 43.720000 ;
      RECT 77.510000 42.640000 79.040000 42.970000 ;
      RECT 53.560000 42.640000 75.710000 43.720000 ;
      RECT 8.560000 42.640000 51.760000 43.720000 ;
      RECT 4.330000 42.640000 6.760000 43.720000 ;
      RECT 1.000000 42.640000 2.530000 42.970000 ;
      RECT 1.000000 41.990000 79.040000 42.640000 ;
      RECT 0.000000 41.140000 80.040000 41.990000 ;
      RECT 0.000000 41.000000 79.040000 41.140000 ;
      RECT 79.310000 39.920000 80.040000 40.160000 ;
      RECT 51.560000 39.920000 77.510000 41.000000 ;
      RECT 6.560000 39.920000 49.760000 41.000000 ;
      RECT 2.530000 39.920000 4.595000 41.000000 ;
      RECT 0.000000 39.920000 0.730000 41.000000 ;
      RECT 0.000000 39.310000 79.040000 39.920000 ;
      RECT 1.000000 38.940000 79.040000 39.310000 ;
      RECT 1.000000 38.330000 80.040000 38.940000 ;
      RECT 0.000000 38.280000 80.040000 38.330000 ;
      RECT 77.510000 38.090000 80.040000 38.280000 ;
      RECT 77.510000 37.200000 79.040000 38.090000 ;
      RECT 53.560000 37.200000 75.710000 38.280000 ;
      RECT 8.560000 37.200000 51.760000 38.280000 ;
      RECT 4.330000 37.200000 6.760000 38.280000 ;
      RECT 0.000000 37.200000 2.530000 38.280000 ;
      RECT 0.000000 37.110000 79.040000 37.200000 ;
      RECT 0.000000 36.870000 80.040000 37.110000 ;
      RECT 0.000000 35.890000 79.040000 36.870000 ;
      RECT 0.000000 35.560000 80.040000 35.890000 ;
      RECT 79.310000 35.040000 80.040000 35.560000 ;
      RECT 0.000000 35.040000 0.730000 35.560000 ;
      RECT 51.560000 34.480000 77.510000 35.560000 ;
      RECT 6.560000 34.480000 49.760000 35.560000 ;
      RECT 2.530000 34.480000 4.595000 35.560000 ;
      RECT 1.000000 34.060000 79.040000 34.480000 ;
      RECT 0.000000 33.820000 80.040000 34.060000 ;
      RECT 0.000000 32.840000 79.040000 33.820000 ;
      RECT 77.510000 31.990000 80.040000 32.840000 ;
      RECT 77.510000 31.760000 79.040000 31.990000 ;
      RECT 53.560000 31.760000 75.710000 32.840000 ;
      RECT 8.560000 31.760000 51.760000 32.840000 ;
      RECT 4.330000 31.760000 6.760000 32.840000 ;
      RECT 0.000000 31.760000 2.530000 32.840000 ;
      RECT 0.000000 31.010000 79.040000 31.760000 ;
      RECT 0.000000 30.770000 80.040000 31.010000 ;
      RECT 1.000000 30.120000 79.040000 30.770000 ;
      RECT 79.310000 29.550000 80.040000 29.790000 ;
      RECT 51.560000 29.040000 77.510000 30.120000 ;
      RECT 6.560000 29.040000 49.760000 30.120000 ;
      RECT 2.530000 29.040000 4.595000 30.120000 ;
      RECT 0.000000 29.040000 0.730000 29.790000 ;
      RECT 0.000000 28.570000 79.040000 29.040000 ;
      RECT 0.000000 27.720000 80.040000 28.570000 ;
      RECT 0.000000 27.400000 79.040000 27.720000 ;
      RECT 77.510000 26.740000 79.040000 27.400000 ;
      RECT 77.510000 26.500000 80.040000 26.740000 ;
      RECT 0.000000 26.500000 2.530000 27.400000 ;
      RECT 77.510000 26.320000 79.040000 26.500000 ;
      RECT 53.560000 26.320000 75.710000 27.400000 ;
      RECT 8.560000 26.320000 51.760000 27.400000 ;
      RECT 4.330000 26.320000 6.760000 27.400000 ;
      RECT 1.000000 26.320000 2.530000 26.500000 ;
      RECT 1.000000 25.520000 79.040000 26.320000 ;
      RECT 0.000000 24.680000 80.040000 25.520000 ;
      RECT 79.310000 24.670000 80.040000 24.680000 ;
      RECT 79.310000 23.600000 80.040000 23.690000 ;
      RECT 51.560000 23.600000 77.510000 24.680000 ;
      RECT 6.560000 23.600000 49.760000 24.680000 ;
      RECT 2.530000 23.600000 4.595000 24.680000 ;
      RECT 0.000000 23.600000 0.730000 24.680000 ;
      RECT 0.000000 23.450000 80.040000 23.600000 ;
      RECT 0.000000 22.470000 79.040000 23.450000 ;
      RECT 0.000000 22.230000 80.040000 22.470000 ;
      RECT 1.000000 21.960000 80.040000 22.230000 ;
      RECT 77.510000 21.620000 80.040000 21.960000 ;
      RECT 1.000000 21.250000 2.530000 21.960000 ;
      RECT 77.510000 20.880000 79.040000 21.620000 ;
      RECT 53.560000 20.880000 75.710000 21.960000 ;
      RECT 8.560000 20.880000 51.760000 21.960000 ;
      RECT 4.330000 20.880000 6.760000 21.960000 ;
      RECT 0.000000 20.880000 2.530000 21.250000 ;
      RECT 0.000000 20.640000 79.040000 20.880000 ;
      RECT 0.000000 20.400000 80.040000 20.640000 ;
      RECT 0.000000 19.420000 79.040000 20.400000 ;
      RECT 0.000000 19.240000 80.040000 19.420000 ;
      RECT 79.310000 18.570000 80.040000 19.240000 ;
      RECT 51.560000 18.160000 77.510000 19.240000 ;
      RECT 6.560000 18.160000 49.760000 19.240000 ;
      RECT 2.530000 18.160000 4.595000 19.240000 ;
      RECT 0.000000 18.160000 0.730000 19.240000 ;
      RECT 0.000000 17.960000 79.040000 18.160000 ;
      RECT 1.000000 17.590000 79.040000 17.960000 ;
      RECT 1.000000 17.350000 80.040000 17.590000 ;
      RECT 1.000000 16.980000 79.040000 17.350000 ;
      RECT 0.000000 16.520000 79.040000 16.980000 ;
      RECT 77.510000 16.370000 79.040000 16.520000 ;
      RECT 77.510000 16.130000 80.040000 16.370000 ;
      RECT 77.510000 15.440000 79.040000 16.130000 ;
      RECT 53.560000 15.440000 75.710000 16.520000 ;
      RECT 8.560000 15.440000 51.760000 16.520000 ;
      RECT 4.330000 15.440000 6.760000 16.520000 ;
      RECT 0.000000 15.440000 2.530000 16.520000 ;
      RECT 0.000000 15.150000 79.040000 15.440000 ;
      RECT 0.000000 14.300000 80.040000 15.150000 ;
      RECT 0.000000 13.800000 79.040000 14.300000 ;
      RECT 0.000000 13.690000 0.730000 13.800000 ;
      RECT 79.310000 13.080000 80.040000 13.320000 ;
      RECT 51.560000 12.720000 77.510000 13.800000 ;
      RECT 6.560000 12.720000 49.760000 13.800000 ;
      RECT 2.530000 12.720000 4.595000 13.800000 ;
      RECT 1.000000 12.710000 79.040000 12.720000 ;
      RECT 0.000000 12.100000 79.040000 12.710000 ;
      RECT 0.000000 11.250000 80.040000 12.100000 ;
      RECT 0.000000 11.080000 79.040000 11.250000 ;
      RECT 77.510000 10.270000 79.040000 11.080000 ;
      RECT 77.510000 10.030000 80.040000 10.270000 ;
      RECT 77.510000 10.000000 79.040000 10.030000 ;
      RECT 53.560000 10.000000 75.710000 11.080000 ;
      RECT 8.560000 10.000000 51.760000 11.080000 ;
      RECT 4.330000 10.000000 6.760000 11.080000 ;
      RECT 0.000000 10.000000 2.530000 11.080000 ;
      RECT 0.000000 9.420000 79.040000 10.000000 ;
      RECT 1.000000 9.050000 79.040000 9.420000 ;
      RECT 1.000000 8.440000 80.040000 9.050000 ;
      RECT 0.000000 8.360000 80.040000 8.440000 ;
      RECT 79.310000 8.200000 80.040000 8.360000 ;
      RECT 51.560000 7.280000 77.510000 8.360000 ;
      RECT 6.560000 7.280000 49.760000 8.360000 ;
      RECT 2.530000 7.280000 4.595000 8.360000 ;
      RECT 0.000000 7.280000 0.730000 8.360000 ;
      RECT 0.000000 7.220000 79.040000 7.280000 ;
      RECT 0.000000 6.980000 80.040000 7.220000 ;
      RECT 0.000000 6.000000 79.040000 6.980000 ;
      RECT 0.000000 5.760000 80.040000 6.000000 ;
      RECT 1.000000 5.640000 79.040000 5.760000 ;
      RECT 77.510000 4.780000 79.040000 5.640000 ;
      RECT 1.000000 4.780000 2.530000 5.640000 ;
      RECT 77.510000 4.560000 80.040000 4.780000 ;
      RECT 53.560000 4.560000 75.710000 5.640000 ;
      RECT 8.560000 4.560000 51.760000 5.640000 ;
      RECT 4.330000 4.560000 6.760000 5.640000 ;
      RECT 0.000000 4.560000 2.530000 4.780000 ;
      RECT 0.000000 4.350000 80.040000 4.560000 ;
      RECT 0.000000 0.000000 80.040000 0.750000 ;
    LAYER met4 ;
      RECT 4.330000 198.320000 75.710000 200.260000 ;
      RECT 51.560000 196.520000 75.710000 198.320000 ;
      RECT 6.560000 196.520000 49.760000 198.320000 ;
      RECT 4.330000 193.320000 4.760000 198.320000 ;
      RECT 4.330000 192.240000 4.595000 193.320000 ;
      RECT 4.330000 187.880000 4.760000 192.240000 ;
      RECT 4.330000 186.800000 4.595000 187.880000 ;
      RECT 4.330000 182.440000 4.760000 186.800000 ;
      RECT 4.330000 181.360000 4.595000 182.440000 ;
      RECT 4.330000 177.000000 4.760000 181.360000 ;
      RECT 4.330000 175.920000 4.595000 177.000000 ;
      RECT 4.330000 171.560000 4.760000 175.920000 ;
      RECT 4.330000 170.480000 4.595000 171.560000 ;
      RECT 4.330000 166.120000 4.760000 170.480000 ;
      RECT 4.330000 165.040000 4.595000 166.120000 ;
      RECT 4.330000 160.680000 4.760000 165.040000 ;
      RECT 4.330000 159.600000 4.595000 160.680000 ;
      RECT 4.330000 155.240000 4.760000 159.600000 ;
      RECT 4.330000 154.160000 4.595000 155.240000 ;
      RECT 4.330000 149.800000 4.760000 154.160000 ;
      RECT 4.330000 148.720000 4.595000 149.800000 ;
      RECT 4.330000 144.360000 4.760000 148.720000 ;
      RECT 4.330000 143.280000 4.595000 144.360000 ;
      RECT 4.330000 138.920000 4.760000 143.280000 ;
      RECT 4.330000 137.840000 4.595000 138.920000 ;
      RECT 4.330000 133.480000 4.760000 137.840000 ;
      RECT 4.330000 132.400000 4.595000 133.480000 ;
      RECT 4.330000 128.040000 4.760000 132.400000 ;
      RECT 4.330000 126.960000 4.595000 128.040000 ;
      RECT 4.330000 122.600000 4.760000 126.960000 ;
      RECT 4.330000 121.520000 4.595000 122.600000 ;
      RECT 4.330000 117.160000 4.760000 121.520000 ;
      RECT 4.330000 116.080000 4.595000 117.160000 ;
      RECT 4.330000 111.720000 4.760000 116.080000 ;
      RECT 4.330000 110.640000 4.595000 111.720000 ;
      RECT 4.330000 106.280000 4.760000 110.640000 ;
      RECT 4.330000 105.200000 4.595000 106.280000 ;
      RECT 4.330000 100.840000 4.760000 105.200000 ;
      RECT 4.330000 99.760000 4.595000 100.840000 ;
      RECT 4.330000 95.400000 4.760000 99.760000 ;
      RECT 4.330000 94.320000 4.595000 95.400000 ;
      RECT 4.330000 89.960000 4.760000 94.320000 ;
      RECT 4.330000 88.880000 4.595000 89.960000 ;
      RECT 4.330000 84.520000 4.760000 88.880000 ;
      RECT 4.330000 83.440000 4.595000 84.520000 ;
      RECT 4.330000 79.080000 4.760000 83.440000 ;
      RECT 4.330000 78.000000 4.595000 79.080000 ;
      RECT 4.330000 73.640000 4.760000 78.000000 ;
      RECT 4.330000 72.560000 4.595000 73.640000 ;
      RECT 4.330000 68.200000 4.760000 72.560000 ;
      RECT 4.330000 67.120000 4.595000 68.200000 ;
      RECT 4.330000 62.760000 4.760000 67.120000 ;
      RECT 4.330000 61.680000 4.595000 62.760000 ;
      RECT 4.330000 57.320000 4.760000 61.680000 ;
      RECT 4.330000 56.240000 4.595000 57.320000 ;
      RECT 4.330000 51.880000 4.760000 56.240000 ;
      RECT 4.330000 50.800000 4.595000 51.880000 ;
      RECT 4.330000 46.440000 4.760000 50.800000 ;
      RECT 4.330000 45.360000 4.595000 46.440000 ;
      RECT 4.330000 41.000000 4.760000 45.360000 ;
      RECT 4.330000 39.920000 4.595000 41.000000 ;
      RECT 4.330000 35.560000 4.760000 39.920000 ;
      RECT 4.330000 34.480000 4.595000 35.560000 ;
      RECT 4.330000 30.120000 4.760000 34.480000 ;
      RECT 4.330000 29.040000 4.595000 30.120000 ;
      RECT 4.330000 24.680000 4.760000 29.040000 ;
      RECT 4.330000 23.600000 4.595000 24.680000 ;
      RECT 4.330000 19.240000 4.760000 23.600000 ;
      RECT 4.330000 18.160000 4.595000 19.240000 ;
      RECT 4.330000 13.800000 4.760000 18.160000 ;
      RECT 4.330000 12.720000 4.595000 13.800000 ;
      RECT 4.330000 8.360000 4.760000 12.720000 ;
      RECT 4.330000 7.280000 4.595000 8.360000 ;
      RECT 53.560000 2.550000 75.710000 196.520000 ;
      RECT 51.560000 2.550000 51.760000 196.520000 ;
      RECT 8.560000 2.550000 49.760000 196.520000 ;
      RECT 6.560000 2.550000 6.760000 196.520000 ;
      RECT 51.560000 0.750000 75.710000 2.550000 ;
      RECT 6.560000 0.750000 49.760000 2.550000 ;
      RECT 4.330000 0.750000 4.760000 7.280000 ;
      RECT 79.310000 0.000000 80.040000 200.260000 ;
      RECT 4.330000 0.000000 75.710000 0.750000 ;
      RECT 0.000000 0.000000 0.730000 200.260000 ;
  END
END W_IO

END LIBRARY
