##
## LEF for PtnCells ;
## created by Innovus v19.11-s128_1 on Wed Nov 24 10:57:13 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO S_term_RAM_IO
  CLASS BLOCK ;
  SIZE 109.940000 BY 30.260000 ;
  FOREIGN S_term_RAM_IO 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6526 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.155 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 8.320000 29.560000 8.700000 30.260000 ;
    END
  END N1BEG[3]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.061 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 6.940000 29.560000 7.320000 30.260000 ;
    END
  END N1BEG[2]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.217 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 6.020000 29.560000 6.400000 30.260000 ;
    END
  END N1BEG[1]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2606 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.195 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 29.560000 5.480000 30.260000 ;
    END
  END N1BEG[0]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.441 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 16.600000 29.560000 16.980000 30.260000 ;
    END
  END N2BEG[7]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 15.680000 29.560000 16.060000 30.260000 ;
    END
  END N2BEG[6]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.313 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 14.760000 29.560000 15.140000 30.260000 ;
    END
  END N2BEG[5]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4966 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.257 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 13.380000 29.560000 13.760000 30.260000 ;
    END
  END N2BEG[4]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6414 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.099 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 12.460000 29.560000 12.840000 30.260000 ;
    END
  END N2BEG[3]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1626 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.705 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 11.540000 29.560000 11.920000 30.260000 ;
    END
  END N2BEG[2]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5602 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.693 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 10.160000 29.560000 10.540000 30.260000 ;
    END
  END N2BEG[1]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2574 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.179 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 9.240000 29.560000 9.620000 30.260000 ;
    END
  END N2BEG[0]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.63 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 25.340000 29.560000 25.720000 30.260000 ;
    END
  END N2BEGb[7]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 24.420000 29.560000 24.800000 30.260000 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.313 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 23.040000 29.560000 23.420000 30.260000 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9982 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.765 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 22.120000 29.560000 22.500000 30.260000 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 21.200000 29.560000 21.580000 30.260000 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7478 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.631 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 19.820000 29.560000 20.200000 30.260000 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.8448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.976 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 18.900000 29.560000 19.280000 30.260000 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.535 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 17.980000 29.560000 18.360000 30.260000 ;
    END
  END N2BEGb[0]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2882 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.333 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 42.820000 29.560000 43.200000 30.260000 ;
    END
  END N4BEG[15]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7478 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.631 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 41.440000 29.560000 41.820000 30.260000 ;
    END
  END N4BEG[14]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5141 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.5678 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.832 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 40.520000 29.560000 40.900000 30.260000 ;
    END
  END N4BEG[13]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7738 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.643 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 39.600000 29.560000 39.980000 30.260000 ;
    END
  END N4BEG[12]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.826 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.904 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 38.220000 29.560000 38.600000 30.260000 ;
    END
  END N4BEG[11]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.077 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.159 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 37.300000 29.560000 37.680000 30.260000 ;
    END
  END N4BEG[10]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0602 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.075 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 36.380000 29.560000 36.760000 30.260000 ;
    END
  END N4BEG[9]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3592 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.678 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 35.000000 29.560000 35.380000 30.260000 ;
    END
  END N4BEG[8]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 29.9316 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 160.576 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 34.080000 29.560000 34.460000 30.260000 ;
    END
  END N4BEG[7]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.313 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 33.160000 29.560000 33.540000 30.260000 ;
    END
  END N4BEG[6]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5362 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.455 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 31.780000 29.560000 32.160000 30.260000 ;
    END
  END N4BEG[5]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6482 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.015 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 30.860000 29.560000 31.240000 30.260000 ;
    END
  END N4BEG[4]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4931 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.024 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 29.940000 29.560000 30.320000 30.260000 ;
    END
  END N4BEG[3]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1725 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.8218 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.52 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 28.560000 29.560000 28.940000 30.260000 ;
    END
  END N4BEG[2]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6849 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.2248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.336 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 27.640000 29.560000 28.020000 30.260000 ;
    END
  END N4BEG[1]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4314 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.049 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 26.260000 29.560000 26.640000 30.260000 ;
    END
  END N4BEG[0]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7384 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.358 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 6.45208 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.741 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.118242 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 46.960000 29.560000 47.340000 30.260000 ;
    END
  END S1END[3]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5838 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.693 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 7.94409 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.1301 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.152078 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 46.040000 29.560000 46.420000 30.260000 ;
    END
  END S1END[2]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.2268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.68 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 15.9846 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 64.8168 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.152221 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 44.660000 29.560000 45.040000 30.260000 ;
    END
  END S1END[1]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8557 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.5568 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.44 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 12.8313 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 48.0375 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203981 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 43.740000 29.560000 44.120000 30.260000 ;
    END
  END S1END[0]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.4522 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.917 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 7.87496 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.3566 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.118242 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 64.440000 29.560000 64.820000 30.260000 ;
    END
  END S2MID[7]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4578 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.063 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 13.9837 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 51.5968 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.170002 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 63.060000 29.560000 63.440000 30.260000 ;
    END
  END S2MID[6]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0602 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.075 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 7.31476 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.5556 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0855958 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 62.140000 29.560000 62.520000 30.260000 ;
    END
  END S2MID[5]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4721 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.9828 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 9.1808 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 45.7614 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.152221 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 61.220000 29.560000 61.600000 30.260000 ;
    END
  END S2MID[4]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7262 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.405 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 16.9098 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 66.2273 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.170002 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 59.840000 29.560000 60.220000 30.260000 ;
    END
  END S2MID[3]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3092 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.342 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 7.10467 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.328 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.6728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.392 LAYER met3  ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 11.0741 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 38.8979 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 58.920000 29.560000 59.300000 30.260000 ;
    END
  END S2MID[2]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7814 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.799 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 9.86405 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.1423 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.152078 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 58.000000 29.560000 58.380000 30.260000 ;
    END
  END S2MID[1]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.205 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 7.23649 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.6093 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.118242 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 56.620000 29.560000 57.000000 30.260000 ;
    END
  END S2MID[0]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 9.39911 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 30.6296 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.119575 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 55.700000 29.560000 56.080000 30.260000 ;
    END
  END S2END[7]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0661 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.1695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.8218 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.52 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 10.3762 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 35.8107 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.152221 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 54.320000 29.560000 54.700000 30.260000 ;
    END
  END S2END[6]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9856 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.702 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 13.614 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 49.7484 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.170002 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 53.400000 29.560000 53.780000 30.260000 ;
    END
  END S2END[5]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.705 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 12.3713 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.4346 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.170002 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 52.480000 29.560000 52.860000 30.260000 ;
    END
  END S2END[4]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2438 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.885 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 6.41007 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.8853 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.118242 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 51.100000 29.560000 51.480000 30.260000 ;
    END
  END S2END[3]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2766 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.039 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 6.02685 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.2783 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.118242 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 50.180000 29.560000 50.560000 30.260000 ;
    END
  END S2END[2]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.535 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 7.41602 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.1621 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0855958 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 49.260000 29.560000 49.640000 30.260000 ;
    END
  END S2END[1]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2982 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.265 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 8.22379 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.8674 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.236485 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 47.880000 29.560000 48.260000 30.260000 ;
    END
  END S2END[0]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3626 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.587 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 8.66133 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.879 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.236485 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 81.460000 29.560000 81.840000 30.260000 ;
    END
  END S4END[15]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5475 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4585 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 8.755 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.0736 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.328502 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.5708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.848 LAYER met3  ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 15.1862 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 59.7729 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.328502 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 80.540000 29.560000 80.920000 30.260000 ;
    END
  END S4END[14]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0674 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.229 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 8.19974 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.0808 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0855958 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 79.620000 29.560000 80.000000 30.260000 ;
    END
  END S4END[13]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0375 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9175 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 7.28548 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.7467 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.328502 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.2808 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.968 LAYER met3  ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 12.6209 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 46.6016 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.328502 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 78.240000 29.560000 78.620000 30.260000 ;
    END
  END S4END[12]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.251 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 7.48737 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.5189 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0855958 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 77.320000 29.560000 77.700000 30.260000 ;
    END
  END S4END[11]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2913 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1775 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 7.72119 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.9045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.328502 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.4308 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.768 LAYER met3  ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 10.6356 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 35.8474 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.328502 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 75.940000 29.560000 76.320000 30.260000 ;
    END
  END S4END[10]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.227 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.027 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 5.59211 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 10.1 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0855958 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 75.020000 29.560000 75.400000 30.260000 ;
    END
  END S4END[9]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.561 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 5.99519 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.3208 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.118242 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 74.100000 29.560000 74.480000 30.260000 ;
    END
  END S4END[8]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.085 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 5.74153 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 10.7897 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0855958 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 72.720000 29.560000 73.100000 30.260000 ;
    END
  END S4END[7]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6006 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.777 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 6.10501 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.1754 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.170002 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 71.800000 29.560000 72.180000 30.260000 ;
    END
  END S4END[6]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.749 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.519 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 8.08752 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.0554 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.236485 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 70.880000 29.560000 71.260000 30.260000 ;
    END
  END S4END[5]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.835 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 7.08583 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.5685 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0855958 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 69.500000 29.560000 69.880000 30.260000 ;
    END
  END S4END[4]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2578 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.955 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 6.01088 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.0211 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.118242 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 68.580000 29.560000 68.960000 30.260000 ;
    END
  END S4END[3]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.691 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.239 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 7.12567 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.5636 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.118242 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 67.660000 29.560000 68.040000 30.260000 ;
    END
  END S4END[2]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0838 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.085 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 7.12363 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.4531 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.118242 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 66.280000 29.560000 66.660000 30.260000 ;
    END
  END S4END[1]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4246 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.907 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 7.56205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.7455 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.118242 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 65.360000 29.560000 65.740000 30.260000 ;
    END
  END S4END[0]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.2416 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.896 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5867 LAYER met3  ;
    ANTENNAMAXAREACAR 9.83101 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 33.6059 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.143452 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 0.000000 5.480000 0.700000 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5724 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.852 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 82.840000 29.560000 83.220000 30.260000 ;
    END
  END UserCLKo
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3458 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.503 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 6.77745 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.5655 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.170002 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 104.460000 0.000000 104.840000 0.700000 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.227 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 6.98999 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 16.8852 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.118242 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 99.400000 0.000000 99.780000 0.700000 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.691 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.239 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 5.79234 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 10.8969 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.118242 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 94.340000 0.000000 94.720000 0.700000 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7482 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.633 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 5.48605 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.94013 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.152078 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 89.280000 0.000000 89.660000 0.700000 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9376 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.462 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 7.9815 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.5858 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.170002 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 84.220000 0.000000 84.600000 0.700000 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5358 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.453 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 10.5258 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.3075 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.170002 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 79.620000 0.000000 80.000000 0.700000 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3996 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.772 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 12.258 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 42.9683 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.170002 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 74.560000 0.000000 74.940000 0.700000 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0598 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.073 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 11.4935 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.1457 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.170002 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 69.500000 0.000000 69.880000 0.700000 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.739 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 8.66058 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.6332 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.170002 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 64.440000 0.000000 64.820000 0.700000 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1074 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.311 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 12.0879 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 42.1176 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.170002 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 59.380000 0.000000 59.760000 0.700000 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.287 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 13.5427 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 49.392 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.170002 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 54.320000 0.000000 54.700000 0.700000 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.6116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.822 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 12.8503 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 45.9215 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.170002 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 49.720000 0.000000 50.100000 0.700000 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3287 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.3645 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 13.6687 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 49.7274 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.2468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.12 LAYER met3  ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 19.8247 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 82.9588 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 44.660000 0.000000 45.040000 0.700000 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9877 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5515 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 8.66552 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.7113 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.7088 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.584 LAYER met3  ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 15.2139 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 60.0358 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 39.600000 0.000000 39.980000 0.700000 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4033 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7375 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 7.43593 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.6565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.5028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.152 LAYER met3  ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 15.5083 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 62.1088 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 34.540000 0.000000 34.920000 0.700000 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5622 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.467 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 6.26946 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.7089 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.118242 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 29.940000 0.000000 30.320000 0.700000 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5622 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.467 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 6.26946 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.3291 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.118242 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 24.880000 0.000000 25.260000 0.700000 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1192 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.1135 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 15.7258 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 59.3892 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.2608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.528 LAYER met3  ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 22.7431 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 97.2146 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 19.820000 0.000000 20.200000 0.700000 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.837 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 20.4206 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 82.5653 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.236485 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 14.760000 0.000000 15.140000 0.700000 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.753 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.421 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 13.9317 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 51.2367 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.170002 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 9.700000 0.000000 10.080000 0.700000 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8902 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 104.460000 29.560000 104.840000 30.260000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 103.080000 29.560000 103.460000 30.260000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4618 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.201 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 102.160000 29.560000 102.540000 30.260000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.271 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.247 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 100.780000 29.560000 101.160000 30.260000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3194 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.489 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.860000 29.560000 100.240000 30.260000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7478 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.631 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 98.940000 29.560000 99.320000 30.260000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.347 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 97.560000 29.560000 97.940000 30.260000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.535 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 96.640000 29.560000 97.020000 30.260000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8218 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.883 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 95.720000 29.560000 96.100000 30.260000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 94.340000 29.560000 94.720000 30.260000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.238 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 93.420000 29.560000 93.800000 30.260000 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0674 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.229 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 92.500000 29.560000 92.880000 30.260000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6526 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.155 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 91.120000 29.560000 91.500000 30.260000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.585 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 90.200000 29.560000 90.580000 30.260000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.371 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 89.280000 29.560000 89.660000 30.260000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.025 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 87.900000 29.560000 88.280000 30.260000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1454 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.619 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 86.980000 29.560000 87.360000 30.260000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3838 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.811 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 86.060000 29.560000 86.440000 30.260000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.019 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.987 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 84.680000 29.560000 85.060000 30.260000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4618 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.201 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 83.760000 29.560000 84.140000 30.260000 ;
    END
  END FrameStrobe_O[0]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 108.740000 25.700000 109.940000 26.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 25.700000 1.200000 26.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.740000 2.850000 109.940000 4.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 1.200000 4.050000 ;
    END
    PORT
      LAYER met4 ;
        RECT 105.910000 29.060000 107.110000 30.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 105.910000 0.000000 107.110000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 29.060000 4.030000 30.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 0.000000 4.030000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 109.940000 4.050000 ;
        RECT 0.000000 25.700000 109.940000 26.900000 ;
        RECT 7.060000 4.860000 8.260000 5.340000 ;
        RECT 2.830000 4.860000 4.030000 5.340000 ;
        RECT 7.060000 10.300000 8.260000 10.780000 ;
        RECT 2.830000 10.300000 4.030000 10.780000 ;
        RECT 52.060000 4.860000 53.260000 5.340000 ;
        RECT 52.060000 10.300000 53.260000 10.780000 ;
        RECT 97.060000 10.300000 98.260000 10.780000 ;
        RECT 97.060000 4.860000 98.260000 5.340000 ;
        RECT 105.910000 10.300000 107.110000 10.780000 ;
        RECT 105.910000 4.860000 107.110000 5.340000 ;
        RECT 7.060000 21.180000 8.260000 21.660000 ;
        RECT 7.060000 15.740000 8.260000 16.220000 ;
        RECT 2.830000 21.180000 4.030000 21.660000 ;
        RECT 2.830000 15.740000 4.030000 16.220000 ;
        RECT 52.060000 15.740000 53.260000 16.220000 ;
        RECT 52.060000 21.180000 53.260000 21.660000 ;
        RECT 97.060000 21.180000 98.260000 21.660000 ;
        RECT 97.060000 15.740000 98.260000 16.220000 ;
        RECT 105.910000 21.180000 107.110000 21.660000 ;
        RECT 105.910000 15.740000 107.110000 16.220000 ;
      LAYER met4 ;
        RECT 97.060000 2.850000 98.260000 26.900000 ;
        RECT 52.060000 2.850000 53.260000 26.900000 ;
        RECT 7.060000 2.850000 8.260000 26.900000 ;
        RECT 105.910000 0.000000 107.110000 30.260000 ;
        RECT 2.830000 0.000000 4.030000 30.260000 ;
    END
# end of P/G power stripe data as pin

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 108.740000 27.500000 109.940000 28.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 27.500000 1.200000 28.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.740000 1.050000 109.940000 2.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 1.200000 2.250000 ;
    END
    PORT
      LAYER met4 ;
        RECT 107.710000 29.060000 108.910000 30.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 107.710000 0.000000 108.910000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 29.060000 2.230000 30.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 0.000000 2.230000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 109.940000 2.250000 ;
        RECT 0.000000 27.500000 109.940000 28.700000 ;
        RECT 1.030000 7.580000 2.230000 8.060000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 1.030000 13.020000 2.230000 13.500000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 50.060000 13.020000 51.260000 13.500000 ;
        RECT 50.060000 7.580000 51.260000 8.060000 ;
        RECT 95.060000 7.580000 96.260000 8.060000 ;
        RECT 95.060000 13.020000 96.260000 13.500000 ;
        RECT 107.710000 7.580000 108.910000 8.060000 ;
        RECT 107.710000 13.020000 108.910000 13.500000 ;
        RECT 1.030000 18.460000 2.230000 18.940000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
        RECT 1.030000 23.900000 2.230000 24.380000 ;
        RECT 50.060000 23.900000 51.260000 24.380000 ;
        RECT 50.060000 18.460000 51.260000 18.940000 ;
        RECT 95.060000 18.460000 96.260000 18.940000 ;
        RECT 95.060000 23.900000 96.260000 24.380000 ;
        RECT 107.710000 18.460000 108.910000 18.940000 ;
        RECT 107.710000 23.900000 108.910000 24.380000 ;
      LAYER met4 ;
        RECT 95.060000 1.050000 96.260000 28.700000 ;
        RECT 50.060000 1.050000 51.260000 28.700000 ;
        RECT 5.060000 1.050000 6.260000 28.700000 ;
        RECT 107.710000 0.000000 108.910000 30.260000 ;
        RECT 1.030000 0.000000 2.230000 30.260000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
    END
# end of P/G power stripe data as pin

  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 109.940000 30.260000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 109.940000 30.260000 ;
    LAYER met2 ;
      RECT 104.980000 29.420000 109.940000 30.260000 ;
      RECT 103.600000 29.420000 104.320000 30.260000 ;
      RECT 102.680000 29.420000 102.940000 30.260000 ;
      RECT 101.300000 29.420000 102.020000 30.260000 ;
      RECT 100.380000 29.420000 100.640000 30.260000 ;
      RECT 99.460000 29.420000 99.720000 30.260000 ;
      RECT 98.080000 29.420000 98.800000 30.260000 ;
      RECT 97.160000 29.420000 97.420000 30.260000 ;
      RECT 96.240000 29.420000 96.500000 30.260000 ;
      RECT 94.860000 29.420000 95.580000 30.260000 ;
      RECT 93.940000 29.420000 94.200000 30.260000 ;
      RECT 93.020000 29.420000 93.280000 30.260000 ;
      RECT 91.640000 29.420000 92.360000 30.260000 ;
      RECT 90.720000 29.420000 90.980000 30.260000 ;
      RECT 89.800000 29.420000 90.060000 30.260000 ;
      RECT 88.420000 29.420000 89.140000 30.260000 ;
      RECT 87.500000 29.420000 87.760000 30.260000 ;
      RECT 86.580000 29.420000 86.840000 30.260000 ;
      RECT 85.200000 29.420000 85.920000 30.260000 ;
      RECT 84.280000 29.420000 84.540000 30.260000 ;
      RECT 83.360000 29.420000 83.620000 30.260000 ;
      RECT 81.980000 29.420000 82.700000 30.260000 ;
      RECT 81.060000 29.420000 81.320000 30.260000 ;
      RECT 80.140000 29.420000 80.400000 30.260000 ;
      RECT 78.760000 29.420000 79.480000 30.260000 ;
      RECT 77.840000 29.420000 78.100000 30.260000 ;
      RECT 76.460000 29.420000 77.180000 30.260000 ;
      RECT 75.540000 29.420000 75.800000 30.260000 ;
      RECT 74.620000 29.420000 74.880000 30.260000 ;
      RECT 73.240000 29.420000 73.960000 30.260000 ;
      RECT 72.320000 29.420000 72.580000 30.260000 ;
      RECT 71.400000 29.420000 71.660000 30.260000 ;
      RECT 70.020000 29.420000 70.740000 30.260000 ;
      RECT 69.100000 29.420000 69.360000 30.260000 ;
      RECT 68.180000 29.420000 68.440000 30.260000 ;
      RECT 66.800000 29.420000 67.520000 30.260000 ;
      RECT 65.880000 29.420000 66.140000 30.260000 ;
      RECT 64.960000 29.420000 65.220000 30.260000 ;
      RECT 63.580000 29.420000 64.300000 30.260000 ;
      RECT 62.660000 29.420000 62.920000 30.260000 ;
      RECT 61.740000 29.420000 62.000000 30.260000 ;
      RECT 60.360000 29.420000 61.080000 30.260000 ;
      RECT 59.440000 29.420000 59.700000 30.260000 ;
      RECT 58.520000 29.420000 58.780000 30.260000 ;
      RECT 57.140000 29.420000 57.860000 30.260000 ;
      RECT 56.220000 29.420000 56.480000 30.260000 ;
      RECT 54.840000 29.420000 55.560000 30.260000 ;
      RECT 53.920000 29.420000 54.180000 30.260000 ;
      RECT 53.000000 29.420000 53.260000 30.260000 ;
      RECT 51.620000 29.420000 52.340000 30.260000 ;
      RECT 50.700000 29.420000 50.960000 30.260000 ;
      RECT 49.780000 29.420000 50.040000 30.260000 ;
      RECT 48.400000 29.420000 49.120000 30.260000 ;
      RECT 47.480000 29.420000 47.740000 30.260000 ;
      RECT 46.560000 29.420000 46.820000 30.260000 ;
      RECT 45.180000 29.420000 45.900000 30.260000 ;
      RECT 44.260000 29.420000 44.520000 30.260000 ;
      RECT 43.340000 29.420000 43.600000 30.260000 ;
      RECT 41.960000 29.420000 42.680000 30.260000 ;
      RECT 41.040000 29.420000 41.300000 30.260000 ;
      RECT 40.120000 29.420000 40.380000 30.260000 ;
      RECT 38.740000 29.420000 39.460000 30.260000 ;
      RECT 37.820000 29.420000 38.080000 30.260000 ;
      RECT 36.900000 29.420000 37.160000 30.260000 ;
      RECT 35.520000 29.420000 36.240000 30.260000 ;
      RECT 34.600000 29.420000 34.860000 30.260000 ;
      RECT 33.680000 29.420000 33.940000 30.260000 ;
      RECT 32.300000 29.420000 33.020000 30.260000 ;
      RECT 31.380000 29.420000 31.640000 30.260000 ;
      RECT 30.460000 29.420000 30.720000 30.260000 ;
      RECT 29.080000 29.420000 29.800000 30.260000 ;
      RECT 28.160000 29.420000 28.420000 30.260000 ;
      RECT 26.780000 29.420000 27.500000 30.260000 ;
      RECT 25.860000 29.420000 26.120000 30.260000 ;
      RECT 24.940000 29.420000 25.200000 30.260000 ;
      RECT 23.560000 29.420000 24.280000 30.260000 ;
      RECT 22.640000 29.420000 22.900000 30.260000 ;
      RECT 21.720000 29.420000 21.980000 30.260000 ;
      RECT 20.340000 29.420000 21.060000 30.260000 ;
      RECT 19.420000 29.420000 19.680000 30.260000 ;
      RECT 18.500000 29.420000 18.760000 30.260000 ;
      RECT 17.120000 29.420000 17.840000 30.260000 ;
      RECT 16.200000 29.420000 16.460000 30.260000 ;
      RECT 15.280000 29.420000 15.540000 30.260000 ;
      RECT 13.900000 29.420000 14.620000 30.260000 ;
      RECT 12.980000 29.420000 13.240000 30.260000 ;
      RECT 12.060000 29.420000 12.320000 30.260000 ;
      RECT 10.680000 29.420000 11.400000 30.260000 ;
      RECT 9.760000 29.420000 10.020000 30.260000 ;
      RECT 8.840000 29.420000 9.100000 30.260000 ;
      RECT 7.460000 29.420000 8.180000 30.260000 ;
      RECT 6.540000 29.420000 6.800000 30.260000 ;
      RECT 5.620000 29.420000 5.880000 30.260000 ;
      RECT 0.000000 29.420000 4.960000 30.260000 ;
      RECT 0.000000 0.840000 109.940000 29.420000 ;
      RECT 104.980000 0.000000 109.940000 0.840000 ;
      RECT 99.920000 0.000000 104.320000 0.840000 ;
      RECT 94.860000 0.000000 99.260000 0.840000 ;
      RECT 89.800000 0.000000 94.200000 0.840000 ;
      RECT 84.740000 0.000000 89.140000 0.840000 ;
      RECT 80.140000 0.000000 84.080000 0.840000 ;
      RECT 75.080000 0.000000 79.480000 0.840000 ;
      RECT 70.020000 0.000000 74.420000 0.840000 ;
      RECT 64.960000 0.000000 69.360000 0.840000 ;
      RECT 59.900000 0.000000 64.300000 0.840000 ;
      RECT 54.840000 0.000000 59.240000 0.840000 ;
      RECT 50.240000 0.000000 54.180000 0.840000 ;
      RECT 45.180000 0.000000 49.580000 0.840000 ;
      RECT 40.120000 0.000000 44.520000 0.840000 ;
      RECT 35.060000 0.000000 39.460000 0.840000 ;
      RECT 30.460000 0.000000 34.400000 0.840000 ;
      RECT 25.400000 0.000000 29.800000 0.840000 ;
      RECT 20.340000 0.000000 24.740000 0.840000 ;
      RECT 15.280000 0.000000 19.680000 0.840000 ;
      RECT 10.220000 0.000000 14.620000 0.840000 ;
      RECT 5.620000 0.000000 9.560000 0.840000 ;
      RECT 0.000000 0.000000 4.960000 0.840000 ;
    LAYER met3 ;
      RECT 0.000000 29.000000 109.940000 30.260000 ;
      RECT 0.000000 24.680000 109.940000 25.400000 ;
      RECT 109.210000 23.600000 109.940000 24.680000 ;
      RECT 96.560000 23.600000 107.410000 24.680000 ;
      RECT 51.560000 23.600000 94.760000 24.680000 ;
      RECT 6.560000 23.600000 49.760000 24.680000 ;
      RECT 2.530000 23.600000 4.595000 24.680000 ;
      RECT 0.000000 23.600000 0.730000 24.680000 ;
      RECT 0.000000 21.960000 109.940000 23.600000 ;
      RECT 107.410000 20.880000 109.940000 21.960000 ;
      RECT 98.560000 20.880000 105.610000 21.960000 ;
      RECT 53.560000 20.880000 96.760000 21.960000 ;
      RECT 8.560000 20.880000 51.760000 21.960000 ;
      RECT 4.330000 20.880000 6.760000 21.960000 ;
      RECT 0.000000 20.880000 2.530000 21.960000 ;
      RECT 0.000000 19.240000 109.940000 20.880000 ;
      RECT 109.210000 18.160000 109.940000 19.240000 ;
      RECT 96.560000 18.160000 107.410000 19.240000 ;
      RECT 51.560000 18.160000 94.760000 19.240000 ;
      RECT 6.560000 18.160000 49.760000 19.240000 ;
      RECT 2.530000 18.160000 4.595000 19.240000 ;
      RECT 0.000000 18.160000 0.730000 19.240000 ;
      RECT 0.000000 16.520000 109.940000 18.160000 ;
      RECT 107.410000 15.440000 109.940000 16.520000 ;
      RECT 98.560000 15.440000 105.610000 16.520000 ;
      RECT 53.560000 15.440000 96.760000 16.520000 ;
      RECT 8.560000 15.440000 51.760000 16.520000 ;
      RECT 4.330000 15.440000 6.760000 16.520000 ;
      RECT 0.000000 15.440000 2.530000 16.520000 ;
      RECT 0.000000 13.800000 109.940000 15.440000 ;
      RECT 109.210000 12.720000 109.940000 13.800000 ;
      RECT 96.560000 12.720000 107.410000 13.800000 ;
      RECT 51.560000 12.720000 94.760000 13.800000 ;
      RECT 6.560000 12.720000 49.760000 13.800000 ;
      RECT 2.530000 12.720000 4.595000 13.800000 ;
      RECT 0.000000 12.720000 0.730000 13.800000 ;
      RECT 0.000000 11.080000 109.940000 12.720000 ;
      RECT 107.410000 10.000000 109.940000 11.080000 ;
      RECT 98.560000 10.000000 105.610000 11.080000 ;
      RECT 53.560000 10.000000 96.760000 11.080000 ;
      RECT 8.560000 10.000000 51.760000 11.080000 ;
      RECT 4.330000 10.000000 6.760000 11.080000 ;
      RECT 0.000000 10.000000 2.530000 11.080000 ;
      RECT 0.000000 8.360000 109.940000 10.000000 ;
      RECT 109.210000 7.280000 109.940000 8.360000 ;
      RECT 96.560000 7.280000 107.410000 8.360000 ;
      RECT 51.560000 7.280000 94.760000 8.360000 ;
      RECT 6.560000 7.280000 49.760000 8.360000 ;
      RECT 2.530000 7.280000 4.595000 8.360000 ;
      RECT 0.000000 7.280000 0.730000 8.360000 ;
      RECT 0.000000 5.640000 109.940000 7.280000 ;
      RECT 107.410000 4.560000 109.940000 5.640000 ;
      RECT 98.560000 4.560000 105.610000 5.640000 ;
      RECT 53.560000 4.560000 96.760000 5.640000 ;
      RECT 8.560000 4.560000 51.760000 5.640000 ;
      RECT 4.330000 4.560000 6.760000 5.640000 ;
      RECT 0.000000 4.560000 2.530000 5.640000 ;
      RECT 0.000000 4.350000 109.940000 4.560000 ;
      RECT 0.000000 0.000000 109.940000 0.750000 ;
    LAYER met4 ;
      RECT 4.330000 29.000000 105.610000 30.260000 ;
      RECT 96.560000 27.200000 105.610000 29.000000 ;
      RECT 51.560000 27.200000 94.760000 29.000000 ;
      RECT 6.560000 27.200000 49.760000 29.000000 ;
      RECT 4.330000 24.680000 4.760000 29.000000 ;
      RECT 4.330000 23.600000 4.595000 24.680000 ;
      RECT 4.330000 19.240000 4.760000 23.600000 ;
      RECT 4.330000 18.160000 4.595000 19.240000 ;
      RECT 4.330000 13.800000 4.760000 18.160000 ;
      RECT 4.330000 12.720000 4.595000 13.800000 ;
      RECT 4.330000 8.360000 4.760000 12.720000 ;
      RECT 4.330000 7.280000 4.595000 8.360000 ;
      RECT 98.560000 2.550000 105.610000 27.200000 ;
      RECT 96.560000 2.550000 96.760000 27.200000 ;
      RECT 53.560000 2.550000 94.760000 27.200000 ;
      RECT 51.560000 2.550000 51.760000 27.200000 ;
      RECT 8.560000 2.550000 49.760000 27.200000 ;
      RECT 6.560000 2.550000 6.760000 27.200000 ;
      RECT 96.560000 0.750000 105.610000 2.550000 ;
      RECT 51.560000 0.750000 94.760000 2.550000 ;
      RECT 6.560000 0.750000 49.760000 2.550000 ;
      RECT 4.330000 0.750000 4.760000 7.280000 ;
      RECT 109.210000 0.000000 109.940000 30.260000 ;
      RECT 4.330000 0.000000 105.610000 0.750000 ;
      RECT 0.000000 0.000000 0.730000 30.260000 ;
  END
END S_term_RAM_IO

END LIBRARY
