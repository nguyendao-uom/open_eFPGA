##
## LEF for PtnCells ;
## created by Innovus v19.11-s128_1 on Tue Nov 23 23:10:52 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO S_term_single2
  CLASS BLOCK ;
  SIZE 200.100000 BY 30.260000 ;
  FOREIGN S_term_single2 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.347 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 9.240000 29.560000 9.620000 30.260000 ;
    END
  END N1BEG[3]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4314 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.049 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 7.860000 29.560000 8.240000 30.260000 ;
    END
  END N1BEG[2]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7455 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.1648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.016 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 6.480000 29.560000 6.860000 30.260000 ;
    END
  END N1BEG[1]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1626 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.705 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 29.560000 5.480000 30.260000 ;
    END
  END N1BEG[0]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1725 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.9508 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.208 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 21.660000 29.560000 22.040000 30.260000 ;
    END
  END N2BEG[7]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7211 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.2928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.032 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 20.280000 29.560000 20.660000 30.260000 ;
    END
  END N2BEG[6]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6526 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.155 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 18.440000 29.560000 18.820000 30.260000 ;
    END
  END N2BEG[5]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1074 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.311 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 17.060000 29.560000 17.440000 30.260000 ;
    END
  END N2BEG[4]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.251 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 15.680000 29.560000 16.060000 30.260000 ;
    END
  END N2BEG[3]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1246 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.397 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 13.840000 29.560000 14.220000 30.260000 ;
    END
  END N2BEG[2]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.441 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 12.460000 29.560000 12.840000 30.260000 ;
    END
  END N2BEG[1]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0602 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.075 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 11.080000 29.560000 11.460000 30.260000 ;
    END
  END N2BEG[0]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.224 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.894 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 34.080000 29.560000 34.460000 30.260000 ;
    END
  END N2BEGb[7]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8694 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.121 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 32.240000 29.560000 32.620000 30.260000 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1288 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.418 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 30.860000 29.560000 31.240000 30.260000 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.553 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 29.480000 29.560000 29.860000 30.260000 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.612 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.952 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 27.640000 29.560000 28.020000 30.260000 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.251 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 26.260000 29.560000 26.640000 30.260000 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.928 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 24.880000 29.560000 25.260000 30.260000 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6849 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.1428 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.232 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 23.040000 29.560000 23.420000 30.260000 ;
    END
  END N2BEGb[0]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2369 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.8258 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.208 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 58.460000 29.560000 58.840000 30.260000 ;
    END
  END N4BEG[15]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.367 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.727 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 56.620000 29.560000 57.000000 30.260000 ;
    END
  END N4BEG[14]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.669 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 55.240000 29.560000 55.620000 30.260000 ;
    END
  END N4BEG[13]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8218 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.883 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 53.860000 29.560000 54.240000 30.260000 ;
    END
  END N4BEG[12]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3458 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.503 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 52.480000 29.560000 52.860000 30.260000 ;
    END
  END N4BEG[11]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.313 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 50.640000 29.560000 51.020000 30.260000 ;
    END
  END N4BEG[10]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8214 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.881 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 49.260000 29.560000 49.640000 30.260000 ;
    END
  END N4BEG[9]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8214 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.881 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 47.880000 29.560000 48.260000 30.260000 ;
    END
  END N4BEG[8]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7455 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.992 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 46.040000 29.560000 46.420000 30.260000 ;
    END
  END N4BEG[7]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7703 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.7548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.496 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 44.660000 29.560000 45.040000 30.260000 ;
    END
  END N4BEG[6]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6954 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.251 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 43.280000 29.560000 43.660000 30.260000 ;
    END
  END N4BEG[5]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7742 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.645 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 41.440000 29.560000 41.820000 30.260000 ;
    END
  END N4BEG[4]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2221 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.9495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.9518 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 90.88 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 40.060000 29.560000 40.440000 30.260000 ;
    END
  END N4BEG[3]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.916 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 38.680000 29.560000 39.060000 30.260000 ;
    END
  END N4BEG[2]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.217 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 36.840000 29.560000 37.220000 30.260000 ;
    END
  END N4BEG[1]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.217 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 35.460000 29.560000 35.840000 30.260000 ;
    END
  END N4BEG[0]
  PIN NN4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0736 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.25 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 82.840000 29.560000 83.220000 30.260000 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.591 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.847 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 81.460000 29.560000 81.840000 30.260000 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.025 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 79.620000 29.560000 80.000000 30.260000 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7262 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.405 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 78.240000 29.560000 78.620000 30.260000 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1762 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.773 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 76.860000 29.560000 77.240000 30.260000 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1246 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.397 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 75.020000 29.560000 75.400000 30.260000 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2842 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.195 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 73.640000 29.560000 74.020000 30.260000 ;
    END
  END NN4BEG[9]
  PIN NN4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0812 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.18 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 72.260000 29.560000 72.640000 30.260000 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1722 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.635 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 70.420000 29.560000 70.800000 30.260000 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0602 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.075 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 69.040000 29.560000 69.420000 30.260000 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6006 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 67.660000 29.560000 68.040000 30.260000 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1343 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.5105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.816 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 65.820000 29.560000 66.200000 30.260000 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4549 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.1135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.7548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.496 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 64.440000 29.560000 64.820000 30.260000 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5838 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.693 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 63.060000 29.560000 63.440000 30.260000 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6395 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.9185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.7098 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.256 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 61.220000 29.560000 61.600000 30.260000 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.665 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.099 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 59.840000 29.560000 60.220000 30.260000 ;
    END
  END NN4BEG[0]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.30626 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.1367 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 88.820000 29.560000 89.200000 30.260000 ;
    END
  END S1END[3]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.313 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.95219 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.31178 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 87.440000 29.560000 87.820000 30.260000 ;
    END
  END S1END[2]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3223 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.5058 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 115.168 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 30.3172 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 160.408 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 86.060000 29.560000 86.440000 30.260000 ;
    END
  END S1END[1]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9807 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.6758 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.408 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 23.2343 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 122.971 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 84.220000 29.560000 84.600000 30.260000 ;
    END
  END S1END[0]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.551 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.15327 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 9.22626 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 113.200000 29.560000 113.580000 30.260000 ;
    END
  END S2MID[7]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3422 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.367 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.06909 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.6465 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 111.820000 29.560000 112.200000 30.260000 ;
    END
  END S2MID[6]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.0128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.872 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 23.5471 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 124.092 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 110.440000 29.560000 110.820000 30.260000 ;
    END
  END S2MID[5]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1058 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.303 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.90721 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 42.996 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 108.600000 29.560000 108.980000 30.260000 ;
    END
  END S2MID[4]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.736 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 11.5397 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 56.3172 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 107.220000 29.560000 107.600000 30.260000 ;
    END
  END S2MID[3]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.9878 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 107.072 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 29.2461 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 153.973 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 105.840000 29.560000 106.220000 30.260000 ;
    END
  END S2MID[2]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9411 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.1108 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 15.9156 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 83.7333 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 104.000000 29.560000 104.380000 30.260000 ;
    END
  END S2MID[1]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7954 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.869 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 11.5095 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 56.1663 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 102.620000 29.560000 103.000000 30.260000 ;
    END
  END S2MID[0]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.157 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.559 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.19583 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.4391 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 101.240000 29.560000 101.620000 30.260000 ;
    END
  END S2END[7]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9959 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.9728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.992 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 17.7076 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 92.6317 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 99.400000 29.560000 99.780000 30.260000 ;
    END
  END S2END[6]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3778 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.663 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.85697 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.7448 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 98.020000 29.560000 98.400000 30.260000 ;
    END
  END S2END[5]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5503 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.3408 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.288 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 21.419 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 113.24 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 96.640000 29.560000 97.020000 30.260000 ;
    END
  END S2END[4]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.371 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.59138 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 36.5758 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 95.260000 29.560000 95.640000 30.260000 ;
    END
  END S2END[3]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8698 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.123 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.82404 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 6.87879 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 93.420000 29.560000 93.800000 30.260000 ;
    END
  END S2END[2]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8694 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.121 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.97791 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.4404 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 92.040000 29.560000 92.420000 30.260000 ;
    END
  END S2END[1]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.145 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.87515 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.08552 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 90.660000 29.560000 91.040000 30.260000 ;
    END
  END S2END[0]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5374 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.461 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.07192 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.8195 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 138.040000 29.560000 138.420000 30.260000 ;
    END
  END S4END[15]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0947 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.3125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.1058 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 118.368 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 32.9278 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 173.731 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 136.200000 29.560000 136.580000 30.260000 ;
    END
  END S4END[14]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3867 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.9858 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 22.2877 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 117.873 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 134.820000 29.560000 135.200000 30.260000 ;
    END
  END S4END[13]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7996 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.89 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.00054 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.6215 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 133.440000 29.560000 133.820000 30.260000 ;
    END
  END S4END[12]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7927 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.4688 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.304 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 15.517 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 81.3845 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 131.600000 29.560000 131.980000 30.260000 ;
    END
  END S4END[11]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2369 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.1908 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.488 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 10.0131 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 51.8532 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 130.220000 29.560000 130.600000 30.260000 ;
    END
  END S4END[10]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7814 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.799 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.7563 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.4067 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 128.840000 29.560000 129.220000 30.260000 ;
    END
  END S4END[9]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1367 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.6428 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 137.232 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 37.9976 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 200.758 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 127.000000 29.560000 127.380000 30.260000 ;
    END
  END S4END[8]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.535 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.20162 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.6269 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 125.620000 29.560000 126.000000 30.260000 ;
    END
  END S4END[7]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.5688 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 6.71084 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 34.4148 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 124.240000 29.560000 124.620000 30.260000 ;
    END
  END S4END[6]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0602 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.075 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.21549 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 9.53737 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 122.400000 29.560000 122.780000 30.260000 ;
    END
  END S4END[5]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.313 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.8 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 12.4599 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 121.020000 29.560000 121.400000 30.260000 ;
    END
  END S4END[4]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8218 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.883 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.9138 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.1199 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 119.640000 29.560000 120.020000 30.260000 ;
    END
  END S4END[3]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.837 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.29717 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.5495 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 117.800000 29.560000 118.180000 30.260000 ;
    END
  END S4END[2]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1402 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.475 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.03623 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 28.732 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 116.420000 29.560000 116.800000 30.260000 ;
    END
  END S4END[1]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.347 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.16229 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.4303 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 115.040000 29.560000 115.420000 30.260000 ;
    END
  END S4END[0]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5686 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.617 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.6804 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.862 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 162.420000 29.560000 162.800000 30.260000 ;
    END
  END SS4END[15]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.717 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.477 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.95906 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.4141 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 160.580000 29.560000 160.960000 30.260000 ;
    END
  END SS4END[14]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.017 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.859 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.8703 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 27.9024 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 159.200000 29.560000 159.580000 30.260000 ;
    END
  END SS4END[13]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.3148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.816 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 9.12054 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 47.0882 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 157.820000 29.560000 158.200000 30.260000 ;
    END
  END SS4END[12]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4287 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.9848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.056 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 13.9615 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 72.5596 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 155.980000 29.560000 156.360000 30.260000 ;
    END
  END SS4END[11]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.441 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.979 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.86222 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 12.771 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 154.600000 29.560000 154.980000 30.260000 ;
    END
  END SS4END[10]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.599 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.74155 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 12.1677 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 153.220000 29.560000 153.600000 30.260000 ;
    END
  END SS4END[9]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.347 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.05556 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.0956 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 151.380000 29.560000 151.760000 30.260000 ;
    END
  END SS4END[8]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.921 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.10646 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.08956 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.000000 29.560000 150.380000 30.260000 ;
    END
  END SS4END[7]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.77 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.0528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.752 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 14.4429 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 72.2465 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 148.620000 29.560000 149.000000 30.260000 ;
    END
  END SS4END[6]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.928 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.12269 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.2323 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 146.780000 29.560000 147.160000 30.260000 ;
    END
  END SS4END[5]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0017 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.7778 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.952 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 21.0762 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 110.734 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 145.400000 29.560000 145.780000 30.260000 ;
    END
  END SS4END[4]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2266 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.025 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.80896 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.3724 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 144.020000 29.560000 144.400000 30.260000 ;
    END
  END SS4END[3]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.305 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.417 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 10.5253 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 51.2451 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 142.640000 29.560000 143.020000 30.260000 ;
    END
  END SS4END[2]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5664 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.714 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.48229 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.0168 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 140.800000 29.560000 141.180000 30.260000 ;
    END
  END SS4END[1]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0814 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.299 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.10303 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.134 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 139.420000 29.560000 139.800000 30.260000 ;
    END
  END SS4END[0]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.152 LAYER met3  ;
    ANTENNAMAXAREACAR 2.16855 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 9.50868 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.0793403 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 0.000000 5.480000 0.700000 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2728 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.354 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 163.800000 29.560000 164.180000 30.260000 ;
    END
  END UserCLKo
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6522 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.153 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.05535 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.8956 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 194.620000 0.000000 195.000000 0.700000 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6074 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.929 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.55946 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.4162 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 184.960000 0.000000 185.340000 0.700000 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6522 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.153 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.83475 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.7926 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 175.300000 0.000000 175.680000 0.700000 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.781 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.797 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.70209 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 27.1293 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 166.100000 0.000000 166.480000 0.700000 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5948 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.866 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.84316 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.1387 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 156.440000 0.000000 156.820000 0.700000 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.781 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.797 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.34559 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.3468 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 147.240000 0.000000 147.620000 0.700000 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8902 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.343 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.39603 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.3077 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 137.580000 0.000000 137.960000 0.700000 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6646 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.097 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.04889 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.7953 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 127.920000 0.000000 128.300000 0.700000 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2632 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.198 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.85508 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.9717 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 118.720000 0.000000 119.100000 0.700000 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0188 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.868 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.61414 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.2276 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 109.060000 0.000000 109.440000 0.700000 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7738 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.643 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.33293 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.1246 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 99.400000 0.000000 99.780000 0.700000 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.525 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.65279 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.7239 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 90.200000 0.000000 90.580000 0.700000 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.1888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.144 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 9.88411 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 47.8559 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 80.540000 0.000000 80.920000 0.700000 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.75 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.524 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.31785 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.0492 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 71.340000 0.000000 71.720000 0.700000 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.869 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.119 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.91178 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.0189 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 61.680000 0.000000 62.060000 0.700000 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7347 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.1048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 139.696 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 38.4117 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 202.945 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 52.480000 0.000000 52.860000 0.700000 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1074 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.311 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.29845 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.0431 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 42.820000 0.000000 43.200000 0.700000 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6931 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.5378 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.672 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 28.5211 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 149.197 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 33.160000 0.000000 33.540000 0.700000 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9678 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.721 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.45724 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.9825 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 23.960000 0.000000 24.340000 0.700000 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5568 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.558 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.9037 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.0694 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 14.300000 0.000000 14.680000 0.700000 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3194 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.489 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 194.160000 29.560000 194.540000 30.260000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6526 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.155 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 192.780000 29.560000 193.160000 30.260000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.367 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.727 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 191.400000 29.560000 191.780000 30.260000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.251 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 190.020000 29.560000 190.400000 30.260000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.717 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.477 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 188.180000 29.560000 188.560000 30.260000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.238 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 186.800000 29.560000 187.180000 30.260000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.217 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 185.420000 29.560000 185.800000 30.260000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0017 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.6728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.392 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 183.580000 29.560000 183.960000 30.260000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.347 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 182.200000 29.560000 182.580000 30.260000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.217 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 180.820000 29.560000 181.200000 30.260000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.217 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 178.980000 29.560000 179.360000 30.260000 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6174 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.861 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 177.600000 29.560000 177.980000 30.260000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.217 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 176.220000 29.560000 176.600000 30.260000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5694 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.621 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 174.380000 29.560000 174.760000 30.260000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.916 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 173.000000 29.560000 173.380000 30.260000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7954 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.869 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 171.620000 29.560000 172.000000 30.260000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8557 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.2488 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.464 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 169.780000 29.560000 170.160000 30.260000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8137 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.9075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.5708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.848 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 168.400000 29.560000 168.780000 30.260000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.553 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 167.020000 29.560000 167.400000 30.260000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.205 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 165.180000 29.560000 165.560000 30.260000 ;
    END
  END FrameStrobe_O[0]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 198.900000 25.700000 200.100000 26.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 25.700000 1.200000 26.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.900000 2.850000 200.100000 4.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 1.200000 4.050000 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.070000 29.060000 197.270000 30.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.070000 0.000000 197.270000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 29.060000 4.030000 30.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 0.000000 4.030000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 200.100000 4.050000 ;
        RECT 0.000000 25.700000 200.100000 26.900000 ;
        RECT 7.060000 4.860000 8.260000 5.340000 ;
        RECT 2.830000 4.860000 4.030000 5.340000 ;
        RECT 7.060000 10.300000 8.260000 10.780000 ;
        RECT 2.830000 10.300000 4.030000 10.780000 ;
        RECT 52.060000 10.300000 53.260000 10.780000 ;
        RECT 97.060000 10.300000 98.260000 10.780000 ;
        RECT 97.060000 4.860000 98.260000 5.340000 ;
        RECT 52.060000 4.860000 53.260000 5.340000 ;
        RECT 142.060000 10.300000 143.260000 10.780000 ;
        RECT 142.060000 4.860000 143.260000 5.340000 ;
        RECT 187.060000 4.860000 188.260000 5.340000 ;
        RECT 187.060000 10.300000 188.260000 10.780000 ;
        RECT 196.070000 10.300000 197.270000 10.780000 ;
        RECT 196.070000 4.860000 197.270000 5.340000 ;
        RECT 2.830000 21.180000 4.030000 21.660000 ;
        RECT 7.060000 21.180000 8.260000 21.660000 ;
        RECT 7.060000 15.740000 8.260000 16.220000 ;
        RECT 2.830000 15.740000 4.030000 16.220000 ;
        RECT 52.060000 21.180000 53.260000 21.660000 ;
        RECT 97.060000 21.180000 98.260000 21.660000 ;
        RECT 97.060000 15.740000 98.260000 16.220000 ;
        RECT 52.060000 15.740000 53.260000 16.220000 ;
        RECT 142.060000 21.180000 143.260000 21.660000 ;
        RECT 142.060000 15.740000 143.260000 16.220000 ;
        RECT 187.060000 15.740000 188.260000 16.220000 ;
        RECT 187.060000 21.180000 188.260000 21.660000 ;
        RECT 196.070000 21.180000 197.270000 21.660000 ;
        RECT 196.070000 15.740000 197.270000 16.220000 ;
      LAYER met4 ;
        RECT 187.060000 2.850000 188.260000 26.900000 ;
        RECT 142.060000 2.850000 143.260000 26.900000 ;
        RECT 97.060000 2.850000 98.260000 26.900000 ;
        RECT 52.060000 2.850000 53.260000 26.900000 ;
        RECT 7.060000 2.850000 8.260000 26.900000 ;
        RECT 196.070000 0.000000 197.270000 30.260000 ;
        RECT 2.830000 0.000000 4.030000 30.260000 ;
    END
# end of P/G power stripe data as pin

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 198.900000 27.500000 200.100000 28.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 27.500000 1.200000 28.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.900000 1.050000 200.100000 2.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 1.200000 2.250000 ;
    END
    PORT
      LAYER met4 ;
        RECT 197.870000 29.060000 199.070000 30.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 197.870000 0.000000 199.070000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 29.060000 2.230000 30.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 0.000000 2.230000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 200.100000 2.250000 ;
        RECT 0.000000 27.500000 200.100000 28.700000 ;
        RECT 1.030000 7.580000 2.230000 8.060000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 1.030000 13.020000 2.230000 13.500000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 50.060000 13.020000 51.260000 13.500000 ;
        RECT 95.060000 13.020000 96.260000 13.500000 ;
        RECT 50.060000 7.580000 51.260000 8.060000 ;
        RECT 95.060000 7.580000 96.260000 8.060000 ;
        RECT 140.060000 13.020000 141.260000 13.500000 ;
        RECT 140.060000 7.580000 141.260000 8.060000 ;
        RECT 185.060000 7.580000 186.260000 8.060000 ;
        RECT 185.060000 13.020000 186.260000 13.500000 ;
        RECT 197.870000 7.580000 199.070000 8.060000 ;
        RECT 197.870000 13.020000 199.070000 13.500000 ;
        RECT 1.030000 18.460000 2.230000 18.940000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 1.030000 23.900000 2.230000 24.380000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
        RECT 50.060000 23.900000 51.260000 24.380000 ;
        RECT 95.060000 23.900000 96.260000 24.380000 ;
        RECT 50.060000 18.460000 51.260000 18.940000 ;
        RECT 95.060000 18.460000 96.260000 18.940000 ;
        RECT 140.060000 23.900000 141.260000 24.380000 ;
        RECT 140.060000 18.460000 141.260000 18.940000 ;
        RECT 185.060000 18.460000 186.260000 18.940000 ;
        RECT 185.060000 23.900000 186.260000 24.380000 ;
        RECT 197.870000 18.460000 199.070000 18.940000 ;
        RECT 197.870000 23.900000 199.070000 24.380000 ;
      LAYER met4 ;
        RECT 185.060000 1.050000 186.260000 28.700000 ;
        RECT 140.060000 1.050000 141.260000 28.700000 ;
        RECT 95.060000 1.050000 96.260000 28.700000 ;
        RECT 50.060000 1.050000 51.260000 28.700000 ;
        RECT 5.060000 1.050000 6.260000 28.700000 ;
        RECT 197.870000 0.000000 199.070000 30.260000 ;
        RECT 1.030000 0.000000 2.230000 30.260000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
    END
# end of P/G power stripe data as pin

  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 200.100000 30.260000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 200.100000 30.260000 ;
    LAYER met2 ;
      RECT 194.680000 29.420000 200.100000 30.260000 ;
      RECT 193.300000 29.420000 194.020000 30.260000 ;
      RECT 191.920000 29.420000 192.640000 30.260000 ;
      RECT 190.540000 29.420000 191.260000 30.260000 ;
      RECT 188.700000 29.420000 189.880000 30.260000 ;
      RECT 187.320000 29.420000 188.040000 30.260000 ;
      RECT 185.940000 29.420000 186.660000 30.260000 ;
      RECT 184.100000 29.420000 185.280000 30.260000 ;
      RECT 182.720000 29.420000 183.440000 30.260000 ;
      RECT 181.340000 29.420000 182.060000 30.260000 ;
      RECT 179.500000 29.420000 180.680000 30.260000 ;
      RECT 178.120000 29.420000 178.840000 30.260000 ;
      RECT 176.740000 29.420000 177.460000 30.260000 ;
      RECT 174.900000 29.420000 176.080000 30.260000 ;
      RECT 173.520000 29.420000 174.240000 30.260000 ;
      RECT 172.140000 29.420000 172.860000 30.260000 ;
      RECT 170.300000 29.420000 171.480000 30.260000 ;
      RECT 168.920000 29.420000 169.640000 30.260000 ;
      RECT 167.540000 29.420000 168.260000 30.260000 ;
      RECT 165.700000 29.420000 166.880000 30.260000 ;
      RECT 164.320000 29.420000 165.040000 30.260000 ;
      RECT 162.940000 29.420000 163.660000 30.260000 ;
      RECT 161.100000 29.420000 162.280000 30.260000 ;
      RECT 159.720000 29.420000 160.440000 30.260000 ;
      RECT 158.340000 29.420000 159.060000 30.260000 ;
      RECT 156.500000 29.420000 157.680000 30.260000 ;
      RECT 155.120000 29.420000 155.840000 30.260000 ;
      RECT 153.740000 29.420000 154.460000 30.260000 ;
      RECT 151.900000 29.420000 153.080000 30.260000 ;
      RECT 150.520000 29.420000 151.240000 30.260000 ;
      RECT 149.140000 29.420000 149.860000 30.260000 ;
      RECT 147.300000 29.420000 148.480000 30.260000 ;
      RECT 145.920000 29.420000 146.640000 30.260000 ;
      RECT 144.540000 29.420000 145.260000 30.260000 ;
      RECT 143.160000 29.420000 143.880000 30.260000 ;
      RECT 141.320000 29.420000 142.500000 30.260000 ;
      RECT 139.940000 29.420000 140.660000 30.260000 ;
      RECT 138.560000 29.420000 139.280000 30.260000 ;
      RECT 136.720000 29.420000 137.900000 30.260000 ;
      RECT 135.340000 29.420000 136.060000 30.260000 ;
      RECT 133.960000 29.420000 134.680000 30.260000 ;
      RECT 132.120000 29.420000 133.300000 30.260000 ;
      RECT 130.740000 29.420000 131.460000 30.260000 ;
      RECT 129.360000 29.420000 130.080000 30.260000 ;
      RECT 127.520000 29.420000 128.700000 30.260000 ;
      RECT 126.140000 29.420000 126.860000 30.260000 ;
      RECT 124.760000 29.420000 125.480000 30.260000 ;
      RECT 122.920000 29.420000 124.100000 30.260000 ;
      RECT 121.540000 29.420000 122.260000 30.260000 ;
      RECT 120.160000 29.420000 120.880000 30.260000 ;
      RECT 118.320000 29.420000 119.500000 30.260000 ;
      RECT 116.940000 29.420000 117.660000 30.260000 ;
      RECT 115.560000 29.420000 116.280000 30.260000 ;
      RECT 113.720000 29.420000 114.900000 30.260000 ;
      RECT 112.340000 29.420000 113.060000 30.260000 ;
      RECT 110.960000 29.420000 111.680000 30.260000 ;
      RECT 109.120000 29.420000 110.300000 30.260000 ;
      RECT 107.740000 29.420000 108.460000 30.260000 ;
      RECT 106.360000 29.420000 107.080000 30.260000 ;
      RECT 104.520000 29.420000 105.700000 30.260000 ;
      RECT 103.140000 29.420000 103.860000 30.260000 ;
      RECT 101.760000 29.420000 102.480000 30.260000 ;
      RECT 99.920000 29.420000 101.100000 30.260000 ;
      RECT 98.540000 29.420000 99.260000 30.260000 ;
      RECT 97.160000 29.420000 97.880000 30.260000 ;
      RECT 95.780000 29.420000 96.500000 30.260000 ;
      RECT 93.940000 29.420000 95.120000 30.260000 ;
      RECT 92.560000 29.420000 93.280000 30.260000 ;
      RECT 91.180000 29.420000 91.900000 30.260000 ;
      RECT 89.340000 29.420000 90.520000 30.260000 ;
      RECT 87.960000 29.420000 88.680000 30.260000 ;
      RECT 86.580000 29.420000 87.300000 30.260000 ;
      RECT 84.740000 29.420000 85.920000 30.260000 ;
      RECT 83.360000 29.420000 84.080000 30.260000 ;
      RECT 81.980000 29.420000 82.700000 30.260000 ;
      RECT 80.140000 29.420000 81.320000 30.260000 ;
      RECT 78.760000 29.420000 79.480000 30.260000 ;
      RECT 77.380000 29.420000 78.100000 30.260000 ;
      RECT 75.540000 29.420000 76.720000 30.260000 ;
      RECT 74.160000 29.420000 74.880000 30.260000 ;
      RECT 72.780000 29.420000 73.500000 30.260000 ;
      RECT 70.940000 29.420000 72.120000 30.260000 ;
      RECT 69.560000 29.420000 70.280000 30.260000 ;
      RECT 68.180000 29.420000 68.900000 30.260000 ;
      RECT 66.340000 29.420000 67.520000 30.260000 ;
      RECT 64.960000 29.420000 65.680000 30.260000 ;
      RECT 63.580000 29.420000 64.300000 30.260000 ;
      RECT 61.740000 29.420000 62.920000 30.260000 ;
      RECT 60.360000 29.420000 61.080000 30.260000 ;
      RECT 58.980000 29.420000 59.700000 30.260000 ;
      RECT 57.140000 29.420000 58.320000 30.260000 ;
      RECT 55.760000 29.420000 56.480000 30.260000 ;
      RECT 54.380000 29.420000 55.100000 30.260000 ;
      RECT 53.000000 29.420000 53.720000 30.260000 ;
      RECT 51.160000 29.420000 52.340000 30.260000 ;
      RECT 49.780000 29.420000 50.500000 30.260000 ;
      RECT 48.400000 29.420000 49.120000 30.260000 ;
      RECT 46.560000 29.420000 47.740000 30.260000 ;
      RECT 45.180000 29.420000 45.900000 30.260000 ;
      RECT 43.800000 29.420000 44.520000 30.260000 ;
      RECT 41.960000 29.420000 43.140000 30.260000 ;
      RECT 40.580000 29.420000 41.300000 30.260000 ;
      RECT 39.200000 29.420000 39.920000 30.260000 ;
      RECT 37.360000 29.420000 38.540000 30.260000 ;
      RECT 35.980000 29.420000 36.700000 30.260000 ;
      RECT 34.600000 29.420000 35.320000 30.260000 ;
      RECT 32.760000 29.420000 33.940000 30.260000 ;
      RECT 31.380000 29.420000 32.100000 30.260000 ;
      RECT 30.000000 29.420000 30.720000 30.260000 ;
      RECT 28.160000 29.420000 29.340000 30.260000 ;
      RECT 26.780000 29.420000 27.500000 30.260000 ;
      RECT 25.400000 29.420000 26.120000 30.260000 ;
      RECT 23.560000 29.420000 24.740000 30.260000 ;
      RECT 22.180000 29.420000 22.900000 30.260000 ;
      RECT 20.800000 29.420000 21.520000 30.260000 ;
      RECT 18.960000 29.420000 20.140000 30.260000 ;
      RECT 17.580000 29.420000 18.300000 30.260000 ;
      RECT 16.200000 29.420000 16.920000 30.260000 ;
      RECT 14.360000 29.420000 15.540000 30.260000 ;
      RECT 12.980000 29.420000 13.700000 30.260000 ;
      RECT 11.600000 29.420000 12.320000 30.260000 ;
      RECT 9.760000 29.420000 10.940000 30.260000 ;
      RECT 8.380000 29.420000 9.100000 30.260000 ;
      RECT 7.000000 29.420000 7.720000 30.260000 ;
      RECT 5.620000 29.420000 6.340000 30.260000 ;
      RECT 0.000000 29.420000 4.960000 30.260000 ;
      RECT 0.000000 0.840000 200.100000 29.420000 ;
      RECT 195.140000 0.000000 200.100000 0.840000 ;
      RECT 185.480000 0.000000 194.480000 0.840000 ;
      RECT 175.820000 0.000000 184.820000 0.840000 ;
      RECT 166.620000 0.000000 175.160000 0.840000 ;
      RECT 156.960000 0.000000 165.960000 0.840000 ;
      RECT 147.760000 0.000000 156.300000 0.840000 ;
      RECT 138.100000 0.000000 147.100000 0.840000 ;
      RECT 128.440000 0.000000 137.440000 0.840000 ;
      RECT 119.240000 0.000000 127.780000 0.840000 ;
      RECT 109.580000 0.000000 118.580000 0.840000 ;
      RECT 99.920000 0.000000 108.920000 0.840000 ;
      RECT 90.720000 0.000000 99.260000 0.840000 ;
      RECT 81.060000 0.000000 90.060000 0.840000 ;
      RECT 71.860000 0.000000 80.400000 0.840000 ;
      RECT 62.200000 0.000000 71.200000 0.840000 ;
      RECT 53.000000 0.000000 61.540000 0.840000 ;
      RECT 43.340000 0.000000 52.340000 0.840000 ;
      RECT 33.680000 0.000000 42.680000 0.840000 ;
      RECT 24.480000 0.000000 33.020000 0.840000 ;
      RECT 14.820000 0.000000 23.820000 0.840000 ;
      RECT 5.620000 0.000000 14.160000 0.840000 ;
      RECT 0.000000 0.000000 4.960000 0.840000 ;
    LAYER met3 ;
      RECT 0.000000 29.000000 200.100000 30.260000 ;
      RECT 0.000000 24.680000 200.100000 25.400000 ;
      RECT 199.370000 23.600000 200.100000 24.680000 ;
      RECT 186.560000 23.600000 197.570000 24.680000 ;
      RECT 141.560000 23.600000 184.760000 24.680000 ;
      RECT 96.560000 23.600000 139.760000 24.680000 ;
      RECT 51.560000 23.600000 94.760000 24.680000 ;
      RECT 6.560000 23.600000 49.760000 24.680000 ;
      RECT 2.530000 23.600000 4.595000 24.680000 ;
      RECT 0.000000 23.600000 0.730000 24.680000 ;
      RECT 0.000000 21.960000 200.100000 23.600000 ;
      RECT 197.570000 20.880000 200.100000 21.960000 ;
      RECT 188.560000 20.880000 195.770000 21.960000 ;
      RECT 143.560000 20.880000 186.760000 21.960000 ;
      RECT 98.560000 20.880000 141.760000 21.960000 ;
      RECT 53.560000 20.880000 96.760000 21.960000 ;
      RECT 8.560000 20.880000 51.760000 21.960000 ;
      RECT 4.330000 20.880000 6.760000 21.960000 ;
      RECT 0.000000 20.880000 2.530000 21.960000 ;
      RECT 0.000000 19.240000 200.100000 20.880000 ;
      RECT 199.370000 18.160000 200.100000 19.240000 ;
      RECT 186.560000 18.160000 197.570000 19.240000 ;
      RECT 141.560000 18.160000 184.760000 19.240000 ;
      RECT 96.560000 18.160000 139.760000 19.240000 ;
      RECT 51.560000 18.160000 94.760000 19.240000 ;
      RECT 6.560000 18.160000 49.760000 19.240000 ;
      RECT 2.530000 18.160000 4.595000 19.240000 ;
      RECT 0.000000 18.160000 0.730000 19.240000 ;
      RECT 0.000000 16.520000 200.100000 18.160000 ;
      RECT 197.570000 15.440000 200.100000 16.520000 ;
      RECT 188.560000 15.440000 195.770000 16.520000 ;
      RECT 143.560000 15.440000 186.760000 16.520000 ;
      RECT 98.560000 15.440000 141.760000 16.520000 ;
      RECT 53.560000 15.440000 96.760000 16.520000 ;
      RECT 8.560000 15.440000 51.760000 16.520000 ;
      RECT 4.330000 15.440000 6.760000 16.520000 ;
      RECT 0.000000 15.440000 2.530000 16.520000 ;
      RECT 0.000000 13.800000 200.100000 15.440000 ;
      RECT 199.370000 12.720000 200.100000 13.800000 ;
      RECT 186.560000 12.720000 197.570000 13.800000 ;
      RECT 141.560000 12.720000 184.760000 13.800000 ;
      RECT 96.560000 12.720000 139.760000 13.800000 ;
      RECT 51.560000 12.720000 94.760000 13.800000 ;
      RECT 6.560000 12.720000 49.760000 13.800000 ;
      RECT 2.530000 12.720000 4.595000 13.800000 ;
      RECT 0.000000 12.720000 0.730000 13.800000 ;
      RECT 0.000000 11.080000 200.100000 12.720000 ;
      RECT 197.570000 10.000000 200.100000 11.080000 ;
      RECT 188.560000 10.000000 195.770000 11.080000 ;
      RECT 143.560000 10.000000 186.760000 11.080000 ;
      RECT 98.560000 10.000000 141.760000 11.080000 ;
      RECT 53.560000 10.000000 96.760000 11.080000 ;
      RECT 8.560000 10.000000 51.760000 11.080000 ;
      RECT 4.330000 10.000000 6.760000 11.080000 ;
      RECT 0.000000 10.000000 2.530000 11.080000 ;
      RECT 0.000000 8.360000 200.100000 10.000000 ;
      RECT 199.370000 7.280000 200.100000 8.360000 ;
      RECT 186.560000 7.280000 197.570000 8.360000 ;
      RECT 141.560000 7.280000 184.760000 8.360000 ;
      RECT 96.560000 7.280000 139.760000 8.360000 ;
      RECT 51.560000 7.280000 94.760000 8.360000 ;
      RECT 6.560000 7.280000 49.760000 8.360000 ;
      RECT 2.530000 7.280000 4.595000 8.360000 ;
      RECT 0.000000 7.280000 0.730000 8.360000 ;
      RECT 0.000000 5.640000 200.100000 7.280000 ;
      RECT 197.570000 4.560000 200.100000 5.640000 ;
      RECT 188.560000 4.560000 195.770000 5.640000 ;
      RECT 143.560000 4.560000 186.760000 5.640000 ;
      RECT 98.560000 4.560000 141.760000 5.640000 ;
      RECT 53.560000 4.560000 96.760000 5.640000 ;
      RECT 8.560000 4.560000 51.760000 5.640000 ;
      RECT 4.330000 4.560000 6.760000 5.640000 ;
      RECT 0.000000 4.560000 2.530000 5.640000 ;
      RECT 0.000000 4.350000 200.100000 4.560000 ;
      RECT 0.000000 0.000000 200.100000 0.750000 ;
    LAYER met4 ;
      RECT 4.330000 29.000000 195.770000 30.260000 ;
      RECT 186.560000 27.200000 195.770000 29.000000 ;
      RECT 141.560000 27.200000 184.760000 29.000000 ;
      RECT 96.560000 27.200000 139.760000 29.000000 ;
      RECT 51.560000 27.200000 94.760000 29.000000 ;
      RECT 6.560000 27.200000 49.760000 29.000000 ;
      RECT 4.330000 24.680000 4.760000 29.000000 ;
      RECT 4.330000 23.600000 4.595000 24.680000 ;
      RECT 4.330000 19.240000 4.760000 23.600000 ;
      RECT 4.330000 18.160000 4.595000 19.240000 ;
      RECT 4.330000 13.800000 4.760000 18.160000 ;
      RECT 4.330000 12.720000 4.595000 13.800000 ;
      RECT 4.330000 8.360000 4.760000 12.720000 ;
      RECT 4.330000 7.280000 4.595000 8.360000 ;
      RECT 188.560000 2.550000 195.770000 27.200000 ;
      RECT 186.560000 2.550000 186.760000 27.200000 ;
      RECT 143.560000 2.550000 184.760000 27.200000 ;
      RECT 141.560000 2.550000 141.760000 27.200000 ;
      RECT 98.560000 2.550000 139.760000 27.200000 ;
      RECT 96.560000 2.550000 96.760000 27.200000 ;
      RECT 53.560000 2.550000 94.760000 27.200000 ;
      RECT 51.560000 2.550000 51.760000 27.200000 ;
      RECT 8.560000 2.550000 49.760000 27.200000 ;
      RECT 6.560000 2.550000 6.760000 27.200000 ;
      RECT 186.560000 0.750000 195.770000 2.550000 ;
      RECT 141.560000 0.750000 184.760000 2.550000 ;
      RECT 96.560000 0.750000 139.760000 2.550000 ;
      RECT 51.560000 0.750000 94.760000 2.550000 ;
      RECT 6.560000 0.750000 49.760000 2.550000 ;
      RECT 4.330000 0.750000 4.760000 7.280000 ;
      RECT 199.370000 0.000000 200.100000 30.260000 ;
      RECT 4.330000 0.000000 195.770000 0.750000 ;
      RECT 0.000000 0.000000 0.730000 30.260000 ;
  END
END S_term_single2

END LIBRARY
