##
## LEF for PtnCells ;
## created by Innovus v19.11-s128_1 on Tue Nov 23 23:00:03 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO N_term_DSP
  CLASS BLOCK ;
  SIZE 200.100000 BY 30.260000 ;
  FOREIGN N_term_DSP 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.585 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.66229 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.2343 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 9.240000 0.000000 9.620000 0.700000 ;
    END
  END N1END[3]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.837 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.23811 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 9.65051 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 7.860000 0.000000 8.240000 0.700000 ;
    END
  END N1END[2]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.736 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.48801 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.363 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 6.480000 0.000000 6.860000 0.700000 ;
    END
  END N1END[1]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.837 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.82397 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.67071 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 0.000000 5.480000 0.700000 ;
    END
  END N1END[0]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.88 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.05677 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.9091 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 21.660000 0.000000 22.040000 0.700000 ;
    END
  END N2MID[7]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0602 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.075 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.99731 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.4465 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 20.280000 0.000000 20.660000 0.700000 ;
    END
  END N2MID[6]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.251 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.53172 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.2774 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 18.440000 0.000000 18.820000 0.700000 ;
    END
  END N2MID[5]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8434 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.109 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 10.4479 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 50.8586 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 17.060000 0.000000 17.440000 0.700000 ;
    END
  END N2MID[4]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.367 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.727 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.28559 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.7556 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 15.680000 0.000000 16.060000 0.700000 ;
    END
  END N2MID[3]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.2948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.376 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 12.2356 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 63.6202 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 13.840000 0.000000 14.220000 0.700000 ;
    END
  END N2MID[2]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6736 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.26 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.04956 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.8667 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 12.460000 0.000000 12.840000 0.700000 ;
    END
  END N2MID[1]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0428 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.096 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.86465 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.01953 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 11.080000 0.000000 11.460000 0.700000 ;
    END
  END N2MID[0]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7213 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.3668 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.76 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 18.863 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 98.8418 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 34.080000 0.000000 34.460000 0.700000 ;
    END
  END N2END[7]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7478 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.631 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.82707 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.7542 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 32.240000 0.000000 32.620000 0.700000 ;
    END
  END N2END[6]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7742 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.645 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.43731 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.6465 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 30.860000 0.000000 31.240000 0.700000 ;
    END
  END N2END[5]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.599 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.26074 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 9.76364 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 29.480000 0.000000 29.860000 0.700000 ;
    END
  END N2END[4]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.784 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.42034 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 45.7205 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 27.640000 0.000000 28.020000 0.700000 ;
    END
  END N2END[3]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.0638 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.144 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 11.1193 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 57.9354 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 26.260000 0.000000 26.640000 0.700000 ;
    END
  END N2END[2]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.4308 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 5.74249 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 29.5111 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 24.880000 0.000000 25.260000 0.700000 ;
    END
  END N2END[1]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4144 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.846 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.1262 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.0909 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 23.040000 0.000000 23.420000 0.700000 ;
    END
  END N2END[0]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.88 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.32209 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.2357 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 58.460000 0.000000 58.840000 0.700000 ;
    END
  END N4END[15]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4746 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.147 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.60013 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 11.4606 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 56.620000 0.000000 57.000000 0.700000 ;
    END
  END N4END[14]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8218 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.883 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.22424 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.5811 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 55.240000 0.000000 55.620000 0.700000 ;
    END
  END N4END[13]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.743 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.489 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.30842 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.002 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 53.860000 0.000000 54.240000 0.700000 ;
    END
  END N4END[12]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9982 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.765 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.41886 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.5542 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 52.480000 0.000000 52.860000 0.700000 ;
    END
  END N4END[11]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9565 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.0868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 7.86498 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 39.8734 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 50.640000 0.000000 51.020000 0.700000 ;
    END
  END N4END[10]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.051 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.80687 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.4943 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 49.260000 0.000000 49.640000 0.700000 ;
    END
  END N4END[9]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9813 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.7455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.9518 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 90.88 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 25.3592 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 133.665 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 47.880000 0.000000 48.260000 0.700000 ;
    END
  END N4END[8]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0629 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.7648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.216 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 12.4939 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 65.7131 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 46.040000 0.000000 46.420000 0.700000 ;
    END
  END N4END[7]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.905 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 12.7671 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 62.4545 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 44.660000 0.000000 45.040000 0.700000 ;
    END
  END N4END[6]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9737 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.4228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.392 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 21.383 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 112.558 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 43.280000 0.000000 43.660000 0.700000 ;
    END
  END N4END[5]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.3288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.224 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 11.1231 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 57.6242 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 41.440000 0.000000 41.820000 0.700000 ;
    END
  END N4END[4]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8406 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.977 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.63273 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.7145 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 40.060000 0.000000 40.440000 0.700000 ;
    END
  END N4END[3]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.837 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.82397 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.67071 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 38.680000 0.000000 39.060000 0.700000 ;
    END
  END N4END[2]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8168 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.976 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.15037 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.3771 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 36.840000 0.000000 37.220000 0.700000 ;
    END
  END N4END[1]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.599 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.75987 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.35017 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 35.460000 0.000000 35.840000 0.700000 ;
    END
  END N4END[0]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4314 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.28047 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 33.73 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 82.840000 0.000000 83.220000 0.700000 ;
    END
  END NN4END[15]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.40222 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.2337 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 81.460000 0.000000 81.840000 0.700000 ;
    END
  END NN4END[14]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.599 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.75987 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.35017 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 79.620000 0.000000 80.000000 0.700000 ;
    END
  END NN4END[13]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1766 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.775 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.4369 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.8034 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 78.240000 0.000000 78.620000 0.700000 ;
    END
  END NN4END[12]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2982 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.265 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.60579 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 11.4889 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 76.860000 0.000000 77.240000 0.700000 ;
    END
  END NN4END[11]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8214 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.881 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.08646 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 28.8923 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 75.020000 0.000000 75.400000 0.700000 ;
    END
  END NN4END[10]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1498 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.523 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.07596 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.83973 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 73.640000 0.000000 74.020000 0.700000 ;
    END
  END NN4END[9]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9722 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.753 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.59758 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.6067 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 72.260000 0.000000 72.640000 0.700000 ;
    END
  END NN4END[8]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.774 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.77791 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.58586 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 70.420000 0.000000 70.800000 0.700000 ;
    END
  END NN4END[7]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.9488 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.864 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 9.18013 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 46.0323 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 69.040000 0.000000 69.420000 0.700000 ;
    END
  END NN4END[6]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9245 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.4058 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.968 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 6.69697 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 33.2835 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 67.660000 0.000000 68.040000 0.700000 ;
    END
  END NN4END[5]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.5695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.1028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 118.352 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 33.0218 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 174.199 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 65.820000 0.000000 66.200000 0.700000 ;
    END
  END NN4END[4]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.3888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 22.9216 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 120.684 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 64.440000 0.000000 64.820000 0.700000 ;
    END
  END NN4END[3]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6511 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.6838 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.784 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 10.7541 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 55.4896 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 63.060000 0.000000 63.440000 0.700000 ;
    END
  END NN4END[2]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.115 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.48983 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 45.9091 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 61.220000 0.000000 61.600000 0.700000 ;
    END
  END NN4END[1]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6187 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.9325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.8508 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.008 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 23.5898 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 124.323 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 59.840000 0.000000 60.220000 0.700000 ;
    END
  END NN4END[0]
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2943 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.1268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.48 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 88.820000 0.000000 89.200000 0.700000 ;
    END
  END S1BEG[3]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.437 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.8258 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.208 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 87.440000 0.000000 87.820000 0.700000 ;
    END
  END S1BEG[2]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1246 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.397 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 86.060000 0.000000 86.440000 0.700000 ;
    END
  END S1BEG[1]
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.5826 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.687 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 84.220000 0.000000 84.600000 0.700000 ;
    END
  END S1BEG[0]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0812 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.18 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 113.200000 0.000000 113.580000 0.700000 ;
    END
  END S2BEG[7]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.535 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.449 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 111.820000 0.000000 112.200000 0.700000 ;
    END
  END S2BEG[6]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.3075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.6748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 110.736 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 110.440000 0.000000 110.820000 0.700000 ;
    END
  END S2BEG[5]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.0442 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.995 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 108.600000 0.000000 108.980000 0.700000 ;
    END
  END S2BEG[4]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.837 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 107.220000 0.000000 107.600000 0.700000 ;
    END
  END S2BEG[3]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.1586 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.567 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 105.840000 0.000000 106.220000 0.700000 ;
    END
  END S2BEG[2]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.727 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.409 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 104.000000 0.000000 104.380000 0.700000 ;
    END
  END S2BEG[1]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9737 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.0538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.424 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 102.620000 0.000000 103.000000 0.700000 ;
    END
  END S2BEG[0]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4861 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.2148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.616 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 101.240000 0.000000 101.620000 0.700000 ;
    END
  END S2BEGb[7]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.6774 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.161 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.400000 0.000000 99.780000 0.700000 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.6028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.352 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 98.020000 0.000000 98.400000 0.700000 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.441 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 96.640000 0.000000 97.020000 0.700000 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.585 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 95.260000 0.000000 95.640000 0.700000 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.5138 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.544 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 93.420000 0.000000 93.800000 0.700000 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.051 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 92.040000 0.000000 92.420000 0.700000 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7266 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.407 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 90.660000 0.000000 91.040000 0.700000 ;
    END
  END S2BEGb[0]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.313 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 138.040000 0.000000 138.420000 0.700000 ;
    END
  END S4BEG[15]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.1425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.2796 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.432 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 136.200000 0.000000 136.580000 0.700000 ;
    END
  END S4BEG[14]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.837 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 134.820000 0.000000 135.200000 0.700000 ;
    END
  END S4BEG[13]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.7664 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.606 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 133.440000 0.000000 133.820000 0.700000 ;
    END
  END S4BEG[12]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2623 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.1505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.7488 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.464 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 131.600000 0.000000 131.980000 0.700000 ;
    END
  END S4BEG[11]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.7088 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.584 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 130.220000 0.000000 130.600000 0.700000 ;
    END
  END S4BEG[10]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0194 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.989 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 128.840000 0.000000 129.220000 0.700000 ;
    END
  END S4BEG[9]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0454 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.001 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 127.000000 0.000000 127.380000 0.700000 ;
    END
  END S4BEG[8]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1445 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.3288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.224 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 125.620000 0.000000 126.000000 0.700000 ;
    END
  END S4BEG[7]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.2468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.12 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 124.240000 0.000000 124.620000 0.700000 ;
    END
  END S4BEG[6]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2092 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.82 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 122.400000 0.000000 122.780000 0.700000 ;
    END
  END S4BEG[5]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.784 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 121.020000 0.000000 121.400000 0.700000 ;
    END
  END S4BEG[4]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.739 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 119.640000 0.000000 120.020000 0.700000 ;
    END
  END S4BEG[3]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8067 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.9388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.144 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 117.800000 0.000000 118.180000 0.700000 ;
    END
  END S4BEG[2]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.298 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 116.420000 0.000000 116.800000 0.700000 ;
    END
  END S4BEG[1]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.217 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 115.040000 0.000000 115.420000 0.700000 ;
    END
  END S4BEG[0]
  PIN SS4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4746 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.147 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 162.420000 0.000000 162.800000 0.700000 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7742 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.645 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 160.580000 0.000000 160.960000 0.700000 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6526 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.155 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 159.200000 0.000000 159.580000 0.700000 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5838 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.693 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.820000 0.000000 158.200000 0.700000 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8434 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.109 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 155.980000 0.000000 156.360000 0.700000 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.605 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.917 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 154.600000 0.000000 154.980000 0.700000 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.837 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 153.220000 0.000000 153.600000 0.700000 ;
    END
  END SS4BEG[9]
  PIN SS4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.536 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 151.380000 0.000000 151.760000 0.700000 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9174 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.361 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.000000 0.000000 150.380000 0.700000 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.347 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 148.620000 0.000000 149.000000 0.700000 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3458 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.503 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 146.780000 0.000000 147.160000 0.700000 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1766 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.775 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 145.400000 0.000000 145.780000 0.700000 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8029 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.2988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.064 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 144.020000 0.000000 144.400000 0.700000 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8698 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.123 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 142.640000 0.000000 143.020000 0.700000 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0598 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.073 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 140.800000 0.000000 141.180000 0.700000 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.3058 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.768 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 139.420000 0.000000 139.800000 0.700000 ;
    END
  END SS4BEG[0]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2299 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.8128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.472 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.152 LAYER met3  ;
    ANTENNAMAXAREACAR 8.2979 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 42.6163 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.0793403 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 163.800000 0.000000 164.180000 0.700000 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3372 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.676 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 29.560000 5.480000 30.260000 ;
    END
  END UserCLKo
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7474 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.629 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.83475 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.7926 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 194.160000 0.000000 194.540000 0.700000 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2714 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.249 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.92424 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 16.9488 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 192.780000 0.000000 193.160000 0.700000 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6522 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.153 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.72034 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.8242 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 191.400000 0.000000 191.780000 0.700000 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7474 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.629 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.43744 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.8061 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 190.020000 0.000000 190.400000 0.700000 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.546 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.77515 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.6397 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 188.180000 0.000000 188.560000 0.700000 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.869 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.119 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.47811 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.8505 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 186.800000 0.000000 187.180000 0.700000 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8732 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.14 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.52458 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.0828 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 185.420000 0.000000 185.800000 0.700000 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6522 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.153 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 10.6456 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 50.8532 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 183.580000 0.000000 183.960000 0.700000 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8214 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.881 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.39704 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.4451 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 182.200000 0.000000 182.580000 0.700000 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.525 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.68276 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.1778 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 180.820000 0.000000 181.200000 0.700000 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8426 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.105 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 14.2354 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 68.3993 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 178.980000 0.000000 179.360000 0.700000 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7738 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.643 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.7666 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.2929 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 177.600000 0.000000 177.980000 0.700000 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6817 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.4208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 20.1469 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 104.58 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 176.220000 0.000000 176.600000 0.700000 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8525 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.1015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.2078 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.912 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 26.9903 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 142.742 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 174.380000 0.000000 174.760000 0.700000 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4045 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.9888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.744 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 23.2003 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 121.005 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 173.000000 0.000000 173.380000 0.700000 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5715 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.4468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.52 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 30.2878 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 159.627 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 171.620000 0.000000 172.000000 0.700000 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9737 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.0238 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.264 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 34.8298 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 183.653 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 169.780000 0.000000 170.160000 0.700000 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.759 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.569 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.28377 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.8788 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 168.400000 0.000000 168.780000 0.700000 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1282 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.533 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 21.203 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 104.634 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 167.020000 0.000000 167.400000 0.700000 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2375 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.0265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.3158 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 151.488 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 39.2767 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 207.063 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 165.180000 0.000000 165.560000 0.700000 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3194 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.489 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 194.620000 29.560000 195.000000 30.260000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.717 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.477 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 184.960000 29.560000 185.340000 30.260000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4622 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.203 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 175.300000 29.560000 175.680000 30.260000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.251 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 166.100000 29.560000 166.480000 30.260000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.251 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 156.440000 29.560000 156.820000 30.260000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.1208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.448 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 147.240000 29.560000 147.620000 30.260000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.217 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 137.580000 29.560000 137.960000 30.260000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.441 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 127.920000 29.560000 128.300000 30.260000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.154 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 118.720000 29.560000 119.100000 30.260000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.217 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 109.060000 29.560000 109.440000 30.260000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.577 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.400000 29.560000 99.780000 30.260000 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.441 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 90.200000 29.560000 90.580000 30.260000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5572 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.56 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 80.540000 29.560000 80.920000 30.260000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.392 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 71.340000 29.560000 71.720000 30.260000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3838 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.811 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 61.680000 29.560000 62.060000 30.260000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5362 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.455 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 52.480000 29.560000 52.860000 30.260000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6174 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.861 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 42.820000 29.560000 43.200000 30.260000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.217 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 33.160000 29.560000 33.540000 30.260000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.823 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 23.960000 29.560000 24.340000 30.260000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.63 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 14.300000 29.560000 14.680000 30.260000 ;
    END
  END FrameStrobe_O[0]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 198.900000 25.700000 200.100000 26.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 25.700000 1.200000 26.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.900000 2.850000 200.100000 4.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 1.200000 4.050000 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.070000 29.060000 197.270000 30.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.070000 0.000000 197.270000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 29.060000 4.030000 30.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 0.000000 4.030000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 200.100000 4.050000 ;
        RECT 0.000000 25.700000 200.100000 26.900000 ;
        RECT 7.060000 4.860000 8.260000 5.340000 ;
        RECT 2.830000 4.860000 4.030000 5.340000 ;
        RECT 7.060000 10.300000 8.260000 10.780000 ;
        RECT 2.830000 10.300000 4.030000 10.780000 ;
        RECT 52.060000 10.300000 53.260000 10.780000 ;
        RECT 97.060000 10.300000 98.260000 10.780000 ;
        RECT 97.060000 4.860000 98.260000 5.340000 ;
        RECT 52.060000 4.860000 53.260000 5.340000 ;
        RECT 142.060000 10.300000 143.260000 10.780000 ;
        RECT 142.060000 4.860000 143.260000 5.340000 ;
        RECT 187.060000 4.860000 188.260000 5.340000 ;
        RECT 187.060000 10.300000 188.260000 10.780000 ;
        RECT 196.070000 10.300000 197.270000 10.780000 ;
        RECT 196.070000 4.860000 197.270000 5.340000 ;
        RECT 2.830000 21.180000 4.030000 21.660000 ;
        RECT 7.060000 21.180000 8.260000 21.660000 ;
        RECT 7.060000 15.740000 8.260000 16.220000 ;
        RECT 2.830000 15.740000 4.030000 16.220000 ;
        RECT 52.060000 21.180000 53.260000 21.660000 ;
        RECT 97.060000 21.180000 98.260000 21.660000 ;
        RECT 97.060000 15.740000 98.260000 16.220000 ;
        RECT 52.060000 15.740000 53.260000 16.220000 ;
        RECT 142.060000 21.180000 143.260000 21.660000 ;
        RECT 142.060000 15.740000 143.260000 16.220000 ;
        RECT 187.060000 15.740000 188.260000 16.220000 ;
        RECT 187.060000 21.180000 188.260000 21.660000 ;
        RECT 196.070000 21.180000 197.270000 21.660000 ;
        RECT 196.070000 15.740000 197.270000 16.220000 ;
      LAYER met4 ;
        RECT 187.060000 2.850000 188.260000 26.900000 ;
        RECT 142.060000 2.850000 143.260000 26.900000 ;
        RECT 97.060000 2.850000 98.260000 26.900000 ;
        RECT 52.060000 2.850000 53.260000 26.900000 ;
        RECT 7.060000 2.850000 8.260000 26.900000 ;
        RECT 196.070000 0.000000 197.270000 30.260000 ;
        RECT 2.830000 0.000000 4.030000 30.260000 ;
    END
# end of P/G power stripe data as pin

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 198.900000 27.500000 200.100000 28.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 27.500000 1.200000 28.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.900000 1.050000 200.100000 2.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 1.200000 2.250000 ;
    END
    PORT
      LAYER met4 ;
        RECT 197.870000 29.060000 199.070000 30.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 197.870000 0.000000 199.070000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 29.060000 2.230000 30.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 0.000000 2.230000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 200.100000 2.250000 ;
        RECT 0.000000 27.500000 200.100000 28.700000 ;
        RECT 1.030000 7.580000 2.230000 8.060000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 1.030000 13.020000 2.230000 13.500000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 50.060000 13.020000 51.260000 13.500000 ;
        RECT 95.060000 13.020000 96.260000 13.500000 ;
        RECT 50.060000 7.580000 51.260000 8.060000 ;
        RECT 95.060000 7.580000 96.260000 8.060000 ;
        RECT 140.060000 13.020000 141.260000 13.500000 ;
        RECT 140.060000 7.580000 141.260000 8.060000 ;
        RECT 185.060000 7.580000 186.260000 8.060000 ;
        RECT 185.060000 13.020000 186.260000 13.500000 ;
        RECT 197.870000 7.580000 199.070000 8.060000 ;
        RECT 197.870000 13.020000 199.070000 13.500000 ;
        RECT 1.030000 18.460000 2.230000 18.940000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 1.030000 23.900000 2.230000 24.380000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
        RECT 50.060000 23.900000 51.260000 24.380000 ;
        RECT 95.060000 23.900000 96.260000 24.380000 ;
        RECT 50.060000 18.460000 51.260000 18.940000 ;
        RECT 95.060000 18.460000 96.260000 18.940000 ;
        RECT 140.060000 23.900000 141.260000 24.380000 ;
        RECT 140.060000 18.460000 141.260000 18.940000 ;
        RECT 185.060000 18.460000 186.260000 18.940000 ;
        RECT 185.060000 23.900000 186.260000 24.380000 ;
        RECT 197.870000 18.460000 199.070000 18.940000 ;
        RECT 197.870000 23.900000 199.070000 24.380000 ;
      LAYER met4 ;
        RECT 185.060000 1.050000 186.260000 28.700000 ;
        RECT 140.060000 1.050000 141.260000 28.700000 ;
        RECT 95.060000 1.050000 96.260000 28.700000 ;
        RECT 50.060000 1.050000 51.260000 28.700000 ;
        RECT 5.060000 1.050000 6.260000 28.700000 ;
        RECT 197.870000 0.000000 199.070000 30.260000 ;
        RECT 1.030000 0.000000 2.230000 30.260000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
    END
# end of P/G power stripe data as pin

  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 200.100000 30.260000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 200.100000 30.260000 ;
    LAYER met2 ;
      RECT 195.140000 29.420000 200.100000 30.260000 ;
      RECT 185.480000 29.420000 194.480000 30.260000 ;
      RECT 175.820000 29.420000 184.820000 30.260000 ;
      RECT 166.620000 29.420000 175.160000 30.260000 ;
      RECT 156.960000 29.420000 165.960000 30.260000 ;
      RECT 147.760000 29.420000 156.300000 30.260000 ;
      RECT 138.100000 29.420000 147.100000 30.260000 ;
      RECT 128.440000 29.420000 137.440000 30.260000 ;
      RECT 119.240000 29.420000 127.780000 30.260000 ;
      RECT 109.580000 29.420000 118.580000 30.260000 ;
      RECT 99.920000 29.420000 108.920000 30.260000 ;
      RECT 90.720000 29.420000 99.260000 30.260000 ;
      RECT 81.060000 29.420000 90.060000 30.260000 ;
      RECT 71.860000 29.420000 80.400000 30.260000 ;
      RECT 62.200000 29.420000 71.200000 30.260000 ;
      RECT 53.000000 29.420000 61.540000 30.260000 ;
      RECT 43.340000 29.420000 52.340000 30.260000 ;
      RECT 33.680000 29.420000 42.680000 30.260000 ;
      RECT 24.480000 29.420000 33.020000 30.260000 ;
      RECT 14.820000 29.420000 23.820000 30.260000 ;
      RECT 5.620000 29.420000 14.160000 30.260000 ;
      RECT 0.000000 29.420000 4.960000 30.260000 ;
      RECT 0.000000 0.840000 200.100000 29.420000 ;
      RECT 194.680000 0.000000 200.100000 0.840000 ;
      RECT 193.300000 0.000000 194.020000 0.840000 ;
      RECT 191.920000 0.000000 192.640000 0.840000 ;
      RECT 190.540000 0.000000 191.260000 0.840000 ;
      RECT 188.700000 0.000000 189.880000 0.840000 ;
      RECT 187.320000 0.000000 188.040000 0.840000 ;
      RECT 185.940000 0.000000 186.660000 0.840000 ;
      RECT 184.100000 0.000000 185.280000 0.840000 ;
      RECT 182.720000 0.000000 183.440000 0.840000 ;
      RECT 181.340000 0.000000 182.060000 0.840000 ;
      RECT 179.500000 0.000000 180.680000 0.840000 ;
      RECT 178.120000 0.000000 178.840000 0.840000 ;
      RECT 176.740000 0.000000 177.460000 0.840000 ;
      RECT 174.900000 0.000000 176.080000 0.840000 ;
      RECT 173.520000 0.000000 174.240000 0.840000 ;
      RECT 172.140000 0.000000 172.860000 0.840000 ;
      RECT 170.300000 0.000000 171.480000 0.840000 ;
      RECT 168.920000 0.000000 169.640000 0.840000 ;
      RECT 167.540000 0.000000 168.260000 0.840000 ;
      RECT 165.700000 0.000000 166.880000 0.840000 ;
      RECT 164.320000 0.000000 165.040000 0.840000 ;
      RECT 162.940000 0.000000 163.660000 0.840000 ;
      RECT 161.100000 0.000000 162.280000 0.840000 ;
      RECT 159.720000 0.000000 160.440000 0.840000 ;
      RECT 158.340000 0.000000 159.060000 0.840000 ;
      RECT 156.500000 0.000000 157.680000 0.840000 ;
      RECT 155.120000 0.000000 155.840000 0.840000 ;
      RECT 153.740000 0.000000 154.460000 0.840000 ;
      RECT 151.900000 0.000000 153.080000 0.840000 ;
      RECT 150.520000 0.000000 151.240000 0.840000 ;
      RECT 149.140000 0.000000 149.860000 0.840000 ;
      RECT 147.300000 0.000000 148.480000 0.840000 ;
      RECT 145.920000 0.000000 146.640000 0.840000 ;
      RECT 144.540000 0.000000 145.260000 0.840000 ;
      RECT 143.160000 0.000000 143.880000 0.840000 ;
      RECT 141.320000 0.000000 142.500000 0.840000 ;
      RECT 139.940000 0.000000 140.660000 0.840000 ;
      RECT 138.560000 0.000000 139.280000 0.840000 ;
      RECT 136.720000 0.000000 137.900000 0.840000 ;
      RECT 135.340000 0.000000 136.060000 0.840000 ;
      RECT 133.960000 0.000000 134.680000 0.840000 ;
      RECT 132.120000 0.000000 133.300000 0.840000 ;
      RECT 130.740000 0.000000 131.460000 0.840000 ;
      RECT 129.360000 0.000000 130.080000 0.840000 ;
      RECT 127.520000 0.000000 128.700000 0.840000 ;
      RECT 126.140000 0.000000 126.860000 0.840000 ;
      RECT 124.760000 0.000000 125.480000 0.840000 ;
      RECT 122.920000 0.000000 124.100000 0.840000 ;
      RECT 121.540000 0.000000 122.260000 0.840000 ;
      RECT 120.160000 0.000000 120.880000 0.840000 ;
      RECT 118.320000 0.000000 119.500000 0.840000 ;
      RECT 116.940000 0.000000 117.660000 0.840000 ;
      RECT 115.560000 0.000000 116.280000 0.840000 ;
      RECT 113.720000 0.000000 114.900000 0.840000 ;
      RECT 112.340000 0.000000 113.060000 0.840000 ;
      RECT 110.960000 0.000000 111.680000 0.840000 ;
      RECT 109.120000 0.000000 110.300000 0.840000 ;
      RECT 107.740000 0.000000 108.460000 0.840000 ;
      RECT 106.360000 0.000000 107.080000 0.840000 ;
      RECT 104.520000 0.000000 105.700000 0.840000 ;
      RECT 103.140000 0.000000 103.860000 0.840000 ;
      RECT 101.760000 0.000000 102.480000 0.840000 ;
      RECT 99.920000 0.000000 101.100000 0.840000 ;
      RECT 98.540000 0.000000 99.260000 0.840000 ;
      RECT 97.160000 0.000000 97.880000 0.840000 ;
      RECT 95.780000 0.000000 96.500000 0.840000 ;
      RECT 93.940000 0.000000 95.120000 0.840000 ;
      RECT 92.560000 0.000000 93.280000 0.840000 ;
      RECT 91.180000 0.000000 91.900000 0.840000 ;
      RECT 89.340000 0.000000 90.520000 0.840000 ;
      RECT 87.960000 0.000000 88.680000 0.840000 ;
      RECT 86.580000 0.000000 87.300000 0.840000 ;
      RECT 84.740000 0.000000 85.920000 0.840000 ;
      RECT 83.360000 0.000000 84.080000 0.840000 ;
      RECT 81.980000 0.000000 82.700000 0.840000 ;
      RECT 80.140000 0.000000 81.320000 0.840000 ;
      RECT 78.760000 0.000000 79.480000 0.840000 ;
      RECT 77.380000 0.000000 78.100000 0.840000 ;
      RECT 75.540000 0.000000 76.720000 0.840000 ;
      RECT 74.160000 0.000000 74.880000 0.840000 ;
      RECT 72.780000 0.000000 73.500000 0.840000 ;
      RECT 70.940000 0.000000 72.120000 0.840000 ;
      RECT 69.560000 0.000000 70.280000 0.840000 ;
      RECT 68.180000 0.000000 68.900000 0.840000 ;
      RECT 66.340000 0.000000 67.520000 0.840000 ;
      RECT 64.960000 0.000000 65.680000 0.840000 ;
      RECT 63.580000 0.000000 64.300000 0.840000 ;
      RECT 61.740000 0.000000 62.920000 0.840000 ;
      RECT 60.360000 0.000000 61.080000 0.840000 ;
      RECT 58.980000 0.000000 59.700000 0.840000 ;
      RECT 57.140000 0.000000 58.320000 0.840000 ;
      RECT 55.760000 0.000000 56.480000 0.840000 ;
      RECT 54.380000 0.000000 55.100000 0.840000 ;
      RECT 53.000000 0.000000 53.720000 0.840000 ;
      RECT 51.160000 0.000000 52.340000 0.840000 ;
      RECT 49.780000 0.000000 50.500000 0.840000 ;
      RECT 48.400000 0.000000 49.120000 0.840000 ;
      RECT 46.560000 0.000000 47.740000 0.840000 ;
      RECT 45.180000 0.000000 45.900000 0.840000 ;
      RECT 43.800000 0.000000 44.520000 0.840000 ;
      RECT 41.960000 0.000000 43.140000 0.840000 ;
      RECT 40.580000 0.000000 41.300000 0.840000 ;
      RECT 39.200000 0.000000 39.920000 0.840000 ;
      RECT 37.360000 0.000000 38.540000 0.840000 ;
      RECT 35.980000 0.000000 36.700000 0.840000 ;
      RECT 34.600000 0.000000 35.320000 0.840000 ;
      RECT 32.760000 0.000000 33.940000 0.840000 ;
      RECT 31.380000 0.000000 32.100000 0.840000 ;
      RECT 30.000000 0.000000 30.720000 0.840000 ;
      RECT 28.160000 0.000000 29.340000 0.840000 ;
      RECT 26.780000 0.000000 27.500000 0.840000 ;
      RECT 25.400000 0.000000 26.120000 0.840000 ;
      RECT 23.560000 0.000000 24.740000 0.840000 ;
      RECT 22.180000 0.000000 22.900000 0.840000 ;
      RECT 20.800000 0.000000 21.520000 0.840000 ;
      RECT 18.960000 0.000000 20.140000 0.840000 ;
      RECT 17.580000 0.000000 18.300000 0.840000 ;
      RECT 16.200000 0.000000 16.920000 0.840000 ;
      RECT 14.360000 0.000000 15.540000 0.840000 ;
      RECT 12.980000 0.000000 13.700000 0.840000 ;
      RECT 11.600000 0.000000 12.320000 0.840000 ;
      RECT 9.760000 0.000000 10.940000 0.840000 ;
      RECT 8.380000 0.000000 9.100000 0.840000 ;
      RECT 7.000000 0.000000 7.720000 0.840000 ;
      RECT 5.620000 0.000000 6.340000 0.840000 ;
      RECT 0.000000 0.000000 4.960000 0.840000 ;
    LAYER met3 ;
      RECT 0.000000 29.000000 200.100000 30.260000 ;
      RECT 0.000000 24.680000 200.100000 25.400000 ;
      RECT 199.370000 23.600000 200.100000 24.680000 ;
      RECT 186.560000 23.600000 197.570000 24.680000 ;
      RECT 141.560000 23.600000 184.760000 24.680000 ;
      RECT 96.560000 23.600000 139.760000 24.680000 ;
      RECT 51.560000 23.600000 94.760000 24.680000 ;
      RECT 6.560000 23.600000 49.760000 24.680000 ;
      RECT 2.530000 23.600000 4.595000 24.680000 ;
      RECT 0.000000 23.600000 0.730000 24.680000 ;
      RECT 0.000000 21.960000 200.100000 23.600000 ;
      RECT 197.570000 20.880000 200.100000 21.960000 ;
      RECT 188.560000 20.880000 195.770000 21.960000 ;
      RECT 143.560000 20.880000 186.760000 21.960000 ;
      RECT 98.560000 20.880000 141.760000 21.960000 ;
      RECT 53.560000 20.880000 96.760000 21.960000 ;
      RECT 8.560000 20.880000 51.760000 21.960000 ;
      RECT 4.330000 20.880000 6.760000 21.960000 ;
      RECT 0.000000 20.880000 2.530000 21.960000 ;
      RECT 0.000000 19.240000 200.100000 20.880000 ;
      RECT 199.370000 18.160000 200.100000 19.240000 ;
      RECT 186.560000 18.160000 197.570000 19.240000 ;
      RECT 141.560000 18.160000 184.760000 19.240000 ;
      RECT 96.560000 18.160000 139.760000 19.240000 ;
      RECT 51.560000 18.160000 94.760000 19.240000 ;
      RECT 6.560000 18.160000 49.760000 19.240000 ;
      RECT 2.530000 18.160000 4.595000 19.240000 ;
      RECT 0.000000 18.160000 0.730000 19.240000 ;
      RECT 0.000000 16.520000 200.100000 18.160000 ;
      RECT 197.570000 15.440000 200.100000 16.520000 ;
      RECT 188.560000 15.440000 195.770000 16.520000 ;
      RECT 143.560000 15.440000 186.760000 16.520000 ;
      RECT 98.560000 15.440000 141.760000 16.520000 ;
      RECT 53.560000 15.440000 96.760000 16.520000 ;
      RECT 8.560000 15.440000 51.760000 16.520000 ;
      RECT 4.330000 15.440000 6.760000 16.520000 ;
      RECT 0.000000 15.440000 2.530000 16.520000 ;
      RECT 0.000000 13.800000 200.100000 15.440000 ;
      RECT 199.370000 12.720000 200.100000 13.800000 ;
      RECT 186.560000 12.720000 197.570000 13.800000 ;
      RECT 141.560000 12.720000 184.760000 13.800000 ;
      RECT 96.560000 12.720000 139.760000 13.800000 ;
      RECT 51.560000 12.720000 94.760000 13.800000 ;
      RECT 6.560000 12.720000 49.760000 13.800000 ;
      RECT 2.530000 12.720000 4.595000 13.800000 ;
      RECT 0.000000 12.720000 0.730000 13.800000 ;
      RECT 0.000000 11.080000 200.100000 12.720000 ;
      RECT 197.570000 10.000000 200.100000 11.080000 ;
      RECT 188.560000 10.000000 195.770000 11.080000 ;
      RECT 143.560000 10.000000 186.760000 11.080000 ;
      RECT 98.560000 10.000000 141.760000 11.080000 ;
      RECT 53.560000 10.000000 96.760000 11.080000 ;
      RECT 8.560000 10.000000 51.760000 11.080000 ;
      RECT 4.330000 10.000000 6.760000 11.080000 ;
      RECT 0.000000 10.000000 2.530000 11.080000 ;
      RECT 0.000000 8.360000 200.100000 10.000000 ;
      RECT 199.370000 7.280000 200.100000 8.360000 ;
      RECT 186.560000 7.280000 197.570000 8.360000 ;
      RECT 141.560000 7.280000 184.760000 8.360000 ;
      RECT 96.560000 7.280000 139.760000 8.360000 ;
      RECT 51.560000 7.280000 94.760000 8.360000 ;
      RECT 6.560000 7.280000 49.760000 8.360000 ;
      RECT 2.530000 7.280000 4.595000 8.360000 ;
      RECT 0.000000 7.280000 0.730000 8.360000 ;
      RECT 0.000000 5.640000 200.100000 7.280000 ;
      RECT 197.570000 4.560000 200.100000 5.640000 ;
      RECT 188.560000 4.560000 195.770000 5.640000 ;
      RECT 143.560000 4.560000 186.760000 5.640000 ;
      RECT 98.560000 4.560000 141.760000 5.640000 ;
      RECT 53.560000 4.560000 96.760000 5.640000 ;
      RECT 8.560000 4.560000 51.760000 5.640000 ;
      RECT 4.330000 4.560000 6.760000 5.640000 ;
      RECT 0.000000 4.560000 2.530000 5.640000 ;
      RECT 0.000000 4.350000 200.100000 4.560000 ;
      RECT 0.000000 0.000000 200.100000 0.750000 ;
    LAYER met4 ;
      RECT 4.330000 29.000000 195.770000 30.260000 ;
      RECT 186.560000 27.200000 195.770000 29.000000 ;
      RECT 141.560000 27.200000 184.760000 29.000000 ;
      RECT 96.560000 27.200000 139.760000 29.000000 ;
      RECT 51.560000 27.200000 94.760000 29.000000 ;
      RECT 6.560000 27.200000 49.760000 29.000000 ;
      RECT 4.330000 24.680000 4.760000 29.000000 ;
      RECT 4.330000 23.600000 4.595000 24.680000 ;
      RECT 4.330000 19.240000 4.760000 23.600000 ;
      RECT 4.330000 18.160000 4.595000 19.240000 ;
      RECT 4.330000 13.800000 4.760000 18.160000 ;
      RECT 4.330000 12.720000 4.595000 13.800000 ;
      RECT 4.330000 8.360000 4.760000 12.720000 ;
      RECT 4.330000 7.280000 4.595000 8.360000 ;
      RECT 188.560000 2.550000 195.770000 27.200000 ;
      RECT 186.560000 2.550000 186.760000 27.200000 ;
      RECT 143.560000 2.550000 184.760000 27.200000 ;
      RECT 141.560000 2.550000 141.760000 27.200000 ;
      RECT 98.560000 2.550000 139.760000 27.200000 ;
      RECT 96.560000 2.550000 96.760000 27.200000 ;
      RECT 53.560000 2.550000 94.760000 27.200000 ;
      RECT 51.560000 2.550000 51.760000 27.200000 ;
      RECT 8.560000 2.550000 49.760000 27.200000 ;
      RECT 6.560000 2.550000 6.760000 27.200000 ;
      RECT 186.560000 0.750000 195.770000 2.550000 ;
      RECT 141.560000 0.750000 184.760000 2.550000 ;
      RECT 96.560000 0.750000 139.760000 2.550000 ;
      RECT 51.560000 0.750000 94.760000 2.550000 ;
      RECT 6.560000 0.750000 49.760000 2.550000 ;
      RECT 4.330000 0.750000 4.760000 7.280000 ;
      RECT 199.370000 0.000000 200.100000 30.260000 ;
      RECT 4.330000 0.000000 195.770000 0.750000 ;
      RECT 0.000000 0.000000 0.730000 30.260000 ;
  END
END N_term_DSP

END LIBRARY
