##
## LEF for PtnCells ;
## created by Innovus v19.11-s128_1 on Mon Dec  6 15:08:48 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO E_CPU_IO
  CLASS BLOCK ;
  SIZE 40.020000 BY 200.260000 ;
  FOREIGN E_CPU_IO 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7296 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.9788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 91.024 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 23.9534 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 107.385 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.1862 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 80.720000 0.700000 81.100000 ;
    END
  END E1END[3]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3396 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.4156 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 109.824 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 27.5574 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 128.781 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 79.500000 0.700000 79.880000 ;
    END
  END E1END[2]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.5868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 16.1528 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 67.2538 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.153554 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 77.670000 0.700000 78.050000 ;
    END
  END E1END[1]
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.3058 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 60.768 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 20.3051 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 78.8821 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.153554 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 76.450000 0.700000 76.830000 ;
    END
  END E1END[0]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 6.80883 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 15.9926 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 92.920000 0.700000 93.300000 ;
    END
  END E2MID[7]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8236 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.0398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 86.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 22.8668 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 102.571 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.1862 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 91.090000 0.700000 91.470000 ;
    END
  END E2MID[6]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.713 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.3798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 66.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 19.3367 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 83.398 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.304443 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 89.870000 0.700000 90.250000 ;
    END
  END E2MID[5]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.392 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 8.25305 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 24.4352 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 88.040000 0.700000 88.420000 ;
    END
  END E2MID[4]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 7.20589 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 18.1044 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 86.820000 0.700000 87.200000 ;
    END
  END E2MID[3]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 5.96945 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 11.9047 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.119575 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 84.990000 0.700000 85.370000 ;
    END
  END E2MID[2]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.401 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.0138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 64.544 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 16.4068 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 68.4934 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.1862 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 83.770000 0.700000 84.150000 ;
    END
  END E2MID[1]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 7.30067 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 19.3559 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 81.940000 0.700000 82.320000 ;
    END
  END E2MID[0]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 6.98597 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 16.9749 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 104.510000 0.700000 104.890000 ;
    END
  END E2END[7]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 10.6811 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 35.1903 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203981 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 103.290000 0.700000 103.670000 ;
    END
  END E2END[6]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0976 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.7337 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 105.712 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 22.0835 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 99.7512 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 101.460000 0.700000 101.840000 ;
    END
  END E2END[5]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2654 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.744 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 8.8415 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 26.8921 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 100.240000 0.700000 100.620000 ;
    END
  END E2END[4]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 6.77893 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 15.9121 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 98.410000 0.700000 98.790000 ;
    END
  END E2END[3]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9016 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.0138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 64.544 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 16.7875 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 71.511 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.1862 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 97.190000 0.700000 97.570000 ;
    END
  END E2END[2]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.9204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.904 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 20.0452 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 55.9628 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.186057 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 95.360000 0.700000 95.740000 ;
    END
  END E2END[1]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 7.00621 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 16.7564 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 94.140000 0.700000 94.520000 ;
    END
  END E2END[0]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 12.8066 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 45.827 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.270464 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 128.300000 0.700000 128.680000 ;
    END
  END EE4END[15]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.088 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 20.7302 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 86.7495 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.2598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 97.856 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 36.2414 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 169.876 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 127.080000 0.700000 127.460000 ;
    END
  END EE4END[14]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.2854 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.984 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 19.5597 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 82.3787 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.0658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 107.488 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 36.6051 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 173.687 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 125.250000 0.700000 125.630000 ;
    END
  END EE4END[13]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.104 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 11.2238 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 38.9326 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.7478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 105.792 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 27.9991 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 128.8 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 124.030000 0.700000 124.410000 ;
    END
  END EE4END[12]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.9584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.44 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 17.2624 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 71.5142 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.152221 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 122.200000 0.700000 122.580000 ;
    END
  END EE4END[11]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6596 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.4518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 50.88 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 18.595 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 78.8526 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.1862 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 120.980000 0.700000 121.360000 ;
    END
  END EE4END[10]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 10.7962 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 36.0331 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.186057 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 119.150000 0.700000 119.530000 ;
    END
  END EE4END[9]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 13.4026 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 48.7447 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203981 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 117.930000 0.700000 118.310000 ;
    END
  END EE4END[8]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 19.6501 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 79.8303 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.42052 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 116.710000 0.700000 117.090000 ;
    END
  END EE4END[7]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 11.5155 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 39.4592 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.152221 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 114.880000 0.700000 115.260000 ;
    END
  END EE4END[6]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 12.6129 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 44.7183 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203981 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 113.660000 0.700000 114.040000 ;
    END
  END EE4END[5]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 12.5927 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 44.7628 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203981 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 111.830000 0.700000 112.210000 ;
    END
  END EE4END[4]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.408 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 9.78797 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 30.9737 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203981 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 110.610000 0.700000 110.990000 ;
    END
  END EE4END[3]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 10.4837 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 34.1725 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203981 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 108.780000 0.700000 109.160000 ;
    END
  END EE4END[2]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 6.60477 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 15.1892 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.119575 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 107.560000 0.700000 107.940000 ;
    END
  END EE4END[1]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.9468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.52 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 16.5814 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 64.658 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 105.730000 0.700000 106.110000 ;
    END
  END EE4END[0]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 18.5954 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 80.7747 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.644758 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 145.990000 0.700000 146.370000 ;
    END
  END E6END[11]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 11.572 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 46.7072 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.466186 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 144.770000 0.700000 145.150000 ;
    END
  END E6END[10]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 11.5335 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 39.7372 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.466186 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 143.550000 0.700000 143.930000 ;
    END
  END E6END[9]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 14.0908 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 58.2708 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.644758 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 141.720000 0.700000 142.100000 ;
    END
  END E6END[8]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.9294 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.952 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 13.0828 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 56.2192 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.466186 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 140.500000 0.700000 140.880000 ;
    END
  END E6END[7]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 13.3552 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 48.0682 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.466186 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 138.670000 0.700000 139.050000 ;
    END
  END E6END[6]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 26.473 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 122.603 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.644758 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 137.450000 0.700000 137.830000 ;
    END
  END E6END[5]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 17.2562 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 67.3803 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.466186 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 135.620000 0.700000 136.000000 ;
    END
  END E6END[4]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.2644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.072 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 20.5566 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 85.1671 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.466186 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 134.400000 0.700000 134.780000 ;
    END
  END E6END[3]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 19.9703 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 89.1833 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.644758 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 132.570000 0.700000 132.950000 ;
    END
  END E6END[2]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.0674 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.688 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 14.3545 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 60.6837 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.466186 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 131.350000 0.700000 131.730000 ;
    END
  END E6END[1]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.5514 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.936 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 31.5274 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 146.882 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.644758 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 130.130000 0.700000 130.510000 ;
    END
  END E6END[0]
  PIN W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.656 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 9.350000 0.700000 9.730000 ;
    END
  END W1BEG[3]
  PIN W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 7.520000 0.700000 7.900000 ;
    END
  END W1BEG[2]
  PIN W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 6.300000 0.700000 6.680000 ;
    END
  END W1BEG[1]
  PIN W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 5.080000 0.700000 5.460000 ;
    END
  END W1BEG[0]
  PIN W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.4834 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 20.940000 0.700000 21.320000 ;
    END
  END W2BEG[7]
  PIN W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 19.720000 0.700000 20.100000 ;
    END
  END W2BEG[6]
  PIN W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.3485 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.096 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 17.890000 0.700000 18.270000 ;
    END
  END W2BEG[5]
  PIN W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.8024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.608 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 16.670000 0.700000 17.050000 ;
    END
  END W2BEG[4]
  PIN W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 15.450000 0.700000 15.830000 ;
    END
  END W2BEG[3]
  PIN W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.3548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.096 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 13.620000 0.700000 14.000000 ;
    END
  END W2BEG[2]
  PIN W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 12.400000 0.700000 12.780000 ;
    END
  END W2BEG[1]
  PIN W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.3114 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.656 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 10.570000 0.700000 10.950000 ;
    END
  END W2BEG[0]
  PIN W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.1964 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.376 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 33.140000 0.700000 33.520000 ;
    END
  END W2BEGb[7]
  PIN W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 31.310000 0.700000 31.690000 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 30.090000 0.700000 30.470000 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.3225 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.576 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 28.870000 0.700000 29.250000 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.3794 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.352 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 27.040000 0.700000 27.420000 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 25.820000 0.700000 26.200000 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 23.990000 0.700000 24.370000 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 22.770000 0.700000 23.150000 ;
    END
  END W2BEGb[0]
  PIN WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 56.930000 0.700000 57.310000 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.6252 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.8 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 55.100000 0.700000 55.480000 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 53.880000 0.700000 54.260000 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.712 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 52.660000 0.700000 53.040000 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 50.830000 0.700000 51.210000 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3046 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.4258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.408 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 49.610000 0.700000 49.990000 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 47.780000 0.700000 48.160000 ;
    END
  END WW4BEG[9]
  PIN WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 46.560000 0.700000 46.940000 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 44.730000 0.700000 45.110000 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 43.510000 0.700000 43.890000 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 42.290000 0.700000 42.670000 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.8384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.8 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 40.460000 0.700000 40.840000 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.0224 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.448 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 39.240000 0.700000 39.620000 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 37.410000 0.700000 37.790000 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 36.190000 0.700000 36.570000 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 34.360000 0.700000 34.740000 ;
    END
  END WW4BEG[0]
  PIN W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 74.620000 0.700000 75.000000 ;
    END
  END W6BEG[11]
  PIN W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 73.400000 0.700000 73.780000 ;
    END
  END W6BEG[10]
  PIN W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 71.570000 0.700000 71.950000 ;
    END
  END W6BEG[9]
  PIN W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 70.350000 0.700000 70.730000 ;
    END
  END W6BEG[8]
  PIN W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 68.520000 0.700000 68.900000 ;
    END
  END W6BEG[7]
  PIN W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 67.300000 0.700000 67.680000 ;
    END
  END W6BEG[6]
  PIN W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 66.080000 0.700000 66.460000 ;
    END
  END W6BEG[5]
  PIN W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 64.250000 0.700000 64.630000 ;
    END
  END W6BEG[4]
  PIN W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.2304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.224 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 63.030000 0.700000 63.410000 ;
    END
  END W6BEG[3]
  PIN W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.3004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.264 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 61.200000 0.700000 61.580000 ;
    END
  END W6BEG[2]
  PIN W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 59.980000 0.700000 60.360000 ;
    END
  END W6BEG[1]
  PIN W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.6804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.624 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 58.150000 0.700000 58.530000 ;
    END
  END W6BEG[0]
  PIN OPA_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 10.8335 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 35.2667 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.466186 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 64.250000 40.020000 64.630000 ;
    END
  END OPA_I0
  PIN OPA_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 8.20758 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 22.4002 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.466186 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 67.910000 40.020000 68.290000 ;
    END
  END OPA_I1
  PIN OPA_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 9.30017 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 30.8062 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.466186 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 71.570000 40.020000 71.950000 ;
    END
  END OPA_I2
  PIN OPA_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 10.252 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 32.5264 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.466186 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 75.230000 40.020000 75.610000 ;
    END
  END OPA_I3
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8029 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.5004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.08 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.8947 LAYER met3  ;
    ANTENNAMAXAREACAR 6.5179 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 30.4502 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 0.000000 5.480000 0.700000 ;
    END
  END UserCLK
  PIN OPB_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7574 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.368 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 10.8282 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 39.4614 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.466186 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 49.000000 40.020000 49.380000 ;
    END
  END OPB_I0
  PIN OPB_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.5854 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.784 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 11.267 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 45.9974 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.466186 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 53.270000 40.020000 53.650000 ;
    END
  END OPB_I1
  PIN OPB_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 13.4814 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 56.7388 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.644758 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 56.930000 40.020000 57.310000 ;
    END
  END OPB_I2
  PIN OPB_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 11.3308 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 46.1324 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.644758 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 60.590000 40.020000 60.970000 ;
    END
  END OPB_I3
  PIN RES0_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.9618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 34.360000 40.020000 34.740000 ;
    END
  END RES0_O0
  PIN RES0_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.9534 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.08 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 38.020000 40.020000 38.400000 ;
    END
  END RES0_O1
  PIN RES0_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9936 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.6518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 121.28 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 41.680000 40.020000 42.060000 ;
    END
  END RES0_O2
  PIN RES0_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.1264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.336 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 45.340000 40.020000 45.720000 ;
    END
  END RES0_O3
  PIN RES1_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.496 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.5448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 163.376 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 19.720000 40.020000 20.100000 ;
    END
  END RES1_O0
  PIN RES1_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2116 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.4228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 157.392 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 23.380000 40.020000 23.760000 ;
    END
  END RES1_O1
  PIN RES1_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 27.040000 40.020000 27.420000 ;
    END
  END RES1_O2
  PIN RES1_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 30.700000 40.020000 31.080000 ;
    END
  END RES1_O3
  PIN RES2_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 5.080000 40.020000 5.460000 ;
    END
  END RES2_O0
  PIN RES2_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3726 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.7478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 105.792 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 8.740000 40.020000 9.120000 ;
    END
  END RES2_O1
  PIN RES2_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 12.400000 40.020000 12.780000 ;
    END
  END RES2_O2
  PIN RES2_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 16.060000 40.020000 16.440000 ;
    END
  END RES2_O3
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 4.5209 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.8898 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.216 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 199.560000 5.480000 200.260000 ;
    END
  END UserCLKo
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3362 LAYER met3  ;
    ANTENNAMAXAREACAR 9.47837 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 38.8028 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.353206 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 194.180000 0.700000 194.560000 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3362 LAYER met3  ;
    ANTENNAMAXAREACAR 9.92417 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 47.9426 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.353206 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 192.350000 0.700000 192.730000 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4766 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.6438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.904 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3362 LAYER met4  ;
    ANTENNAMAXAREACAR 18.283 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 89.6473 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.383142 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 191.130000 0.700000 191.510000 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3362 LAYER met3  ;
    ANTENNAMAXAREACAR 9.89739 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 46.9288 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.353206 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 189.300000 0.700000 189.680000 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3362 LAYER met3  ;
    ANTENNAMAXAREACAR 8.848 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 26.4034 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.228535 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 188.080000 0.700000 188.460000 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3362 LAYER met3  ;
    ANTENNAMAXAREACAR 10.9987 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 37.0643 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.353206 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 186.250000 0.700000 186.630000 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3362 LAYER met3  ;
    ANTENNAMAXAREACAR 13.8406 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 50.8404 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.353206 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 185.030000 0.700000 185.410000 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3362 LAYER met3  ;
    ANTENNAMAXAREACAR 11.2556 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 38.2751 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.353206 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 183.200000 0.700000 183.580000 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3362 LAYER met3  ;
    ANTENNAMAXAREACAR 18.7653 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 75.3848 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.353206 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 181.980000 0.700000 182.360000 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3362 LAYER met3  ;
    ANTENNAMAXAREACAR 13.3946 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 63.3775 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.353206 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 180.760000 0.700000 181.140000 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3362 LAYER met3  ;
    ANTENNAMAXAREACAR 10.3849 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 33.9812 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.228535 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 178.930000 0.700000 179.310000 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.8892 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3362 LAYER met3  ;
    ANTENNAMAXAREACAR 15.3513 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 75.209 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 177.710000 0.700000 178.090000 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3362 LAYER met3  ;
    ANTENNAMAXAREACAR 16.6736 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 78.2455 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 175.880000 0.700000 176.260000 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.2836 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.8926 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 144.368 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3362 LAYER met4  ;
    ANTENNAMAXAREACAR 28.6179 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 152.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.458019 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 174.660000 0.700000 175.040000 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6866 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.7727 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 153.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3362 LAYER met4  ;
    ANTENNAMAXAREACAR 30.2325 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 141.424 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.354407 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 172.830000 0.700000 173.210000 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8044 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.752 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 18.143 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 92.5502 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.230842 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.3208 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 92.848 LAYER met4  ;
    ANTENNAGATEAREA 1.3362 LAYER met4  ;
    ANTENNAMAXAREACAR 31.1058 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 162.037 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.458019 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 171.610000 0.700000 171.990000 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7186 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.6698 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 41.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3362 LAYER met4  ;
    ANTENNAMAXAREACAR 17.9529 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 79.568 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.383142 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 169.780000 0.700000 170.160000 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3362 LAYER met3  ;
    ANTENNAMAXAREACAR 11.8404 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 57.6368 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.353206 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 168.560000 0.700000 168.940000 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.2946 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.0407 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 134.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3362 LAYER met4  ;
    ANTENNAMAXAREACAR 30.7289 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 144.592 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.458019 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 167.340000 0.700000 167.720000 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.367 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.0378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 64.672 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3362 LAYER met4  ;
    ANTENNAMAXAREACAR 18.3828 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 83.823 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.383142 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 165.510000 0.700000 165.890000 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 7.48361 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 27.7447 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.152221 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 164.290000 0.700000 164.670000 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 13.9176 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 51.4119 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.270464 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 162.460000 0.700000 162.840000 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.4892 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.408 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 21.3343 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 90.5424 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 161.240000 0.700000 161.620000 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 16.0324 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 61.857 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.270464 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 159.410000 0.700000 159.790000 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 15.9554 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 61.4019 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203981 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 158.190000 0.700000 158.570000 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 11.1601 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 37.2814 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203981 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 156.360000 0.700000 156.740000 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.3188 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 71.504 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 19.8737 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 85.7721 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.23796 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 155.140000 0.700000 155.520000 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.229 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.9528 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 69.552 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 19.2492 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 85.0634 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.23796 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 153.920000 0.700000 154.300000 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1546 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.0748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.536 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 20.0298 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 98.1438 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.1862 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 152.090000 0.700000 152.470000 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.5686 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.024 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.8808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 85.168 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 19.4785 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 89.7345 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.1862 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 150.870000 0.700000 151.250000 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 13.2217 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 47.6811 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203981 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 149.040000 0.700000 149.420000 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3396 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.5888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 88.944 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 20.1084 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 98.6551 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.1862 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 147.820000 0.700000 148.200000 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 193.570000 40.020000 193.950000 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 189.910000 40.020000 190.290000 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 186.250000 40.020000 186.630000 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 182.590000 40.020000 182.970000 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 178.930000 40.020000 179.310000 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 175.270000 40.020000 175.650000 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.9544 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.752 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 171.610000 40.020000 171.990000 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 167.950000 40.020000 168.330000 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 164.290000 40.020000 164.670000 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.7914 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.216 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 160.630000 40.020000 161.010000 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 156.970000 40.020000 157.350000 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 153.310000 40.020000 153.690000 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 149.650000 40.020000 150.030000 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 145.380000 40.020000 145.760000 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 141.720000 40.020000 142.100000 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 138.060000 40.020000 138.440000 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 134.400000 40.020000 134.780000 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 130.740000 40.020000 131.120000 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 127.080000 40.020000 127.460000 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 123.420000 40.020000 123.800000 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.5368 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 119.760000 40.020000 120.140000 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 116.100000 40.020000 116.480000 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 112.440000 40.020000 112.820000 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.664 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 108.780000 40.020000 109.160000 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 105.120000 40.020000 105.500000 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 101.460000 40.020000 101.840000 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 97.190000 40.020000 97.570000 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 93.530000 40.020000 93.910000 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 89.870000 40.020000 90.250000 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 86.210000 40.020000 86.590000 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 82.550000 40.020000 82.930000 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 39.320000 78.890000 40.020000 79.270000 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 19.711 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 98.329 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 23.0851 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 97.1039 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.170002 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 34.540000 0.000000 34.920000 0.700000 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.357 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 121.569 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 25.6391 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 110.131 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.118242 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 32.700000 0.000000 33.080000 0.700000 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1112 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.33 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 8.63102 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.1055 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0855958 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 31.320000 0.000000 31.700000 0.700000 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.1967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.7145 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 16.3106 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.0527 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 17.5482 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 70.7269 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.3936 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 131.04 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 38.2699 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 182.042 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 29.940000 0.000000 30.320000 0.700000 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8454 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.119 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 8.93819 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.7675 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.152078 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 28.560000 0.000000 28.940000 0.700000 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6069 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6965 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 8.49689 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.8256 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 12.1155 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 44.1983 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.4418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 248.16 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 51.5666 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 255.004 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 27.180000 0.000000 27.560000 0.700000 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.879 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.207 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 6.82241 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.7983 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 9.48861 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 31.0916 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.4288 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 253.424 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 49.7781 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 246.368 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 25.340000 0.000000 25.720000 0.700000 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3179 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.3205 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 12.4329 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.6646 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 13.0196 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 47.8238 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.2788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 204.624 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 45.5364 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 221.646 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 23.960000 0.000000 24.340000 0.700000 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.2414 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.981 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 29.8197 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 130.847 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.236485 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 22.580000 0.000000 22.960000 0.700000 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8887 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.1645 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 12.0713 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.7403 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 13.1502 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 48.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.6598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 238.656 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 51.0875 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 251.3 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 21.200000 0.000000 21.580000 0.700000 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.7851 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 83.6465 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 45.4743 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 208.6 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 49.4104 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 230.666 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8568 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 101.04 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 65.4287 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 316.497 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 19.360000 0.000000 19.740000 0.700000 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.3478 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 121.513 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 30.4705 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 134.101 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.236485 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 17.980000 0.000000 18.360000 0.700000 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0277 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.8695 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 16.726 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 65.13 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 19.2335 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 79.5767 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.6098 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 233.056 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 56.2789 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 277.552 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 16.600000 0.000000 16.980000 0.700000 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.129 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.537 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 9.51974 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.6752 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.152078 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 15.220000 0.000000 15.600000 0.700000 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0485 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 9.64987 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.977 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 11.9986 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 43.5772 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.0148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 251.216 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 51.9364 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 256.978 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 13.840000 0.000000 14.220000 0.700000 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7175 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.992 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met3  ;
    ANTENNAMAXAREACAR 10.5185 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 35.3353 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.119575 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 12.460000 0.000000 12.840000 0.700000 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.0458 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 115.003 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1772 LAYER met2  ;
    ANTENNAMAXAREACAR 27.8765 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 121.131 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.236485 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 10.620000 0.000000 11.000000 0.700000 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2661 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0515 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 9.57902 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.1235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 10.1562 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 33.2827 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.2698 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 268.576 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 52.8591 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 261.431 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 9.240000 0.000000 9.620000 0.700000 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5815 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 7.8836 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.5567 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 8.46078 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 24.7159 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.5508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 259.408 LAYER met4  ;
    ANTENNAGATEAREA 1.1772 LAYER met4  ;
    ANTENNAMAXAREACAR 49.7034 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 245.076 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 7.860000 0.000000 8.240000 0.700000 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.0886 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 140.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8112 LAYER met4  ;
    ANTENNAMAXAREACAR 31.9333 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 152.492 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.868344 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 6.480000 0.000000 6.860000 0.700000 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8454 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.119 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 34.540000 199.560000 34.920000 200.260000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.2706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.245 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 32.700000 199.560000 33.080000 200.260000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4989 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.3335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8088 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.784 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 31.320000 199.560000 31.700000 200.260000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8434 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.109 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 29.940000 199.560000 30.320000 200.260000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.3846 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.815 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 28.560000 199.560000 28.940000 200.260000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.6038 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.911 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 27.180000 199.560000 27.560000 200.260000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.8768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 25.340000 199.560000 25.720000 200.260000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.3814 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.799 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 23.960000 199.560000 24.340000 200.260000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.4138 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.961 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 22.580000 199.560000 22.960000 200.260000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7326 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.555 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 21.200000 199.560000 21.580000 200.260000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2738 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.261 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 19.360000 199.560000 19.740000 200.260000 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.4638 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.211 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 17.980000 199.560000 18.360000 200.260000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.9296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.53 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 16.600000 199.560000 16.980000 200.260000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.685 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.317 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 15.220000 199.560000 15.600000 200.260000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.2398 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.091 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 13.840000 199.560000 14.220000 200.260000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.9066 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 12.460000 199.560000 12.840000 200.260000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.4942 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.363 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 10.620000 199.560000 11.000000 200.260000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.2874 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.329 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 9.240000 199.560000 9.620000 200.260000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.3878 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.831 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 7.860000 199.560000 8.240000 200.260000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5574 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.679 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 6.480000 199.560000 6.860000 200.260000 ;
    END
  END FrameStrobe_O[0]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 38.820000 195.020000 40.020000 196.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 195.020000 1.200000 196.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.820000 2.850000 40.020000 4.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 1.200000 4.050000 ;
    END
    PORT
      LAYER met4 ;
        RECT 35.990000 199.060000 37.190000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 35.990000 0.000000 37.190000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 199.060000 4.030000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 0.000000 4.030000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 40.020000 4.050000 ;
        RECT 0.000000 195.020000 40.020000 196.220000 ;
        RECT 2.830000 4.860000 4.030000 5.340000 ;
        RECT 2.830000 10.300000 4.030000 10.780000 ;
        RECT 7.060000 4.860000 8.260000 5.340000 ;
        RECT 7.060000 10.300000 8.260000 10.780000 ;
        RECT 7.060000 21.180000 8.260000 21.660000 ;
        RECT 7.060000 15.740000 8.260000 16.220000 ;
        RECT 2.830000 15.740000 4.030000 16.220000 ;
        RECT 2.830000 21.180000 4.030000 21.660000 ;
        RECT 2.830000 37.500000 4.030000 37.980000 ;
        RECT 7.060000 37.500000 8.260000 37.980000 ;
        RECT 7.060000 32.060000 8.260000 32.540000 ;
        RECT 7.060000 26.620000 8.260000 27.100000 ;
        RECT 2.830000 32.060000 4.030000 32.540000 ;
        RECT 2.830000 26.620000 4.030000 27.100000 ;
        RECT 7.060000 42.940000 8.260000 43.420000 ;
        RECT 7.060000 48.380000 8.260000 48.860000 ;
        RECT 2.830000 48.380000 4.030000 48.860000 ;
        RECT 2.830000 42.940000 4.030000 43.420000 ;
        RECT 7.060000 59.260000 8.260000 59.740000 ;
        RECT 7.060000 53.820000 8.260000 54.300000 ;
        RECT 2.830000 53.820000 4.030000 54.300000 ;
        RECT 2.830000 59.260000 4.030000 59.740000 ;
        RECT 7.060000 70.140000 8.260000 70.620000 ;
        RECT 7.060000 64.700000 8.260000 65.180000 ;
        RECT 2.830000 70.140000 4.030000 70.620000 ;
        RECT 2.830000 64.700000 4.030000 65.180000 ;
        RECT 7.060000 86.460000 8.260000 86.940000 ;
        RECT 7.060000 81.020000 8.260000 81.500000 ;
        RECT 7.060000 75.580000 8.260000 76.060000 ;
        RECT 2.830000 86.460000 4.030000 86.940000 ;
        RECT 2.830000 81.020000 4.030000 81.500000 ;
        RECT 2.830000 75.580000 4.030000 76.060000 ;
        RECT 7.060000 97.340000 8.260000 97.820000 ;
        RECT 7.060000 91.900000 8.260000 92.380000 ;
        RECT 2.830000 97.340000 4.030000 97.820000 ;
        RECT 2.830000 91.900000 4.030000 92.380000 ;
        RECT 35.990000 4.860000 37.190000 5.340000 ;
        RECT 35.990000 10.300000 37.190000 10.780000 ;
        RECT 35.990000 15.740000 37.190000 16.220000 ;
        RECT 35.990000 21.180000 37.190000 21.660000 ;
        RECT 35.990000 37.500000 37.190000 37.980000 ;
        RECT 35.990000 26.620000 37.190000 27.100000 ;
        RECT 35.990000 32.060000 37.190000 32.540000 ;
        RECT 35.990000 42.940000 37.190000 43.420000 ;
        RECT 35.990000 48.380000 37.190000 48.860000 ;
        RECT 35.990000 53.820000 37.190000 54.300000 ;
        RECT 35.990000 59.260000 37.190000 59.740000 ;
        RECT 35.990000 70.140000 37.190000 70.620000 ;
        RECT 35.990000 64.700000 37.190000 65.180000 ;
        RECT 35.990000 86.460000 37.190000 86.940000 ;
        RECT 35.990000 81.020000 37.190000 81.500000 ;
        RECT 35.990000 75.580000 37.190000 76.060000 ;
        RECT 35.990000 97.340000 37.190000 97.820000 ;
        RECT 35.990000 91.900000 37.190000 92.380000 ;
        RECT 7.060000 108.220000 8.260000 108.700000 ;
        RECT 7.060000 102.780000 8.260000 103.260000 ;
        RECT 2.830000 108.220000 4.030000 108.700000 ;
        RECT 2.830000 102.780000 4.030000 103.260000 ;
        RECT 7.060000 124.540000 8.260000 125.020000 ;
        RECT 7.060000 119.100000 8.260000 119.580000 ;
        RECT 7.060000 113.660000 8.260000 114.140000 ;
        RECT 2.830000 124.540000 4.030000 125.020000 ;
        RECT 2.830000 119.100000 4.030000 119.580000 ;
        RECT 2.830000 113.660000 4.030000 114.140000 ;
        RECT 7.060000 129.980000 8.260000 130.460000 ;
        RECT 7.060000 135.420000 8.260000 135.900000 ;
        RECT 2.830000 135.420000 4.030000 135.900000 ;
        RECT 2.830000 129.980000 4.030000 130.460000 ;
        RECT 7.060000 140.860000 8.260000 141.340000 ;
        RECT 7.060000 146.300000 8.260000 146.780000 ;
        RECT 2.830000 140.860000 4.030000 141.340000 ;
        RECT 2.830000 146.300000 4.030000 146.780000 ;
        RECT 2.830000 162.620000 4.030000 163.100000 ;
        RECT 7.060000 162.620000 8.260000 163.100000 ;
        RECT 7.060000 157.180000 8.260000 157.660000 ;
        RECT 7.060000 151.740000 8.260000 152.220000 ;
        RECT 2.830000 157.180000 4.030000 157.660000 ;
        RECT 2.830000 151.740000 4.030000 152.220000 ;
        RECT 7.060000 173.500000 8.260000 173.980000 ;
        RECT 7.060000 168.060000 8.260000 168.540000 ;
        RECT 2.830000 173.500000 4.030000 173.980000 ;
        RECT 2.830000 168.060000 4.030000 168.540000 ;
        RECT 7.060000 184.380000 8.260000 184.860000 ;
        RECT 7.060000 178.940000 8.260000 179.420000 ;
        RECT 2.830000 178.940000 4.030000 179.420000 ;
        RECT 2.830000 184.380000 4.030000 184.860000 ;
        RECT 2.830000 189.820000 4.030000 190.300000 ;
        RECT 7.060000 189.820000 8.260000 190.300000 ;
        RECT 35.990000 102.780000 37.190000 103.260000 ;
        RECT 35.990000 108.220000 37.190000 108.700000 ;
        RECT 35.990000 113.660000 37.190000 114.140000 ;
        RECT 35.990000 119.100000 37.190000 119.580000 ;
        RECT 35.990000 124.540000 37.190000 125.020000 ;
        RECT 35.990000 129.980000 37.190000 130.460000 ;
        RECT 35.990000 135.420000 37.190000 135.900000 ;
        RECT 35.990000 140.860000 37.190000 141.340000 ;
        RECT 35.990000 146.300000 37.190000 146.780000 ;
        RECT 35.990000 162.620000 37.190000 163.100000 ;
        RECT 35.990000 157.180000 37.190000 157.660000 ;
        RECT 35.990000 151.740000 37.190000 152.220000 ;
        RECT 35.990000 173.500000 37.190000 173.980000 ;
        RECT 35.990000 168.060000 37.190000 168.540000 ;
        RECT 35.990000 178.940000 37.190000 179.420000 ;
        RECT 35.990000 184.380000 37.190000 184.860000 ;
        RECT 35.990000 189.820000 37.190000 190.300000 ;
      LAYER met4 ;
        RECT 7.060000 2.850000 8.260000 196.220000 ;
        RECT 35.990000 0.000000 37.190000 200.260000 ;
        RECT 2.830000 0.000000 4.030000 200.260000 ;
    END
# end of P/G power stripe data as pin

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 38.820000 196.820000 40.020000 198.020000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 196.820000 1.200000 198.020000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.820000 1.050000 40.020000 2.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 1.200000 2.250000 ;
    END
    PORT
      LAYER met4 ;
        RECT 37.790000 199.060000 38.990000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 37.790000 0.000000 38.990000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 199.060000 2.230000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 0.000000 2.230000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 40.020000 2.250000 ;
        RECT 0.000000 196.820000 40.020000 198.020000 ;
        RECT 37.790000 100.060000 38.990000 100.540000 ;
        RECT 4.895000 100.060000 6.260000 100.540000 ;
        RECT 1.030000 100.060000 2.230000 100.540000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 1.030000 7.580000 2.230000 8.060000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 1.030000 18.460000 2.230000 18.940000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 1.030000 13.020000 2.230000 13.500000 ;
        RECT 1.030000 23.900000 2.230000 24.380000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
        RECT 1.030000 29.340000 2.230000 29.820000 ;
        RECT 4.895000 29.340000 6.260000 29.820000 ;
        RECT 1.030000 34.780000 2.230000 35.260000 ;
        RECT 4.895000 34.780000 6.260000 35.260000 ;
        RECT 1.030000 40.220000 2.230000 40.700000 ;
        RECT 4.895000 40.220000 6.260000 40.700000 ;
        RECT 1.030000 45.660000 2.230000 46.140000 ;
        RECT 4.895000 45.660000 6.260000 46.140000 ;
        RECT 4.895000 51.100000 6.260000 51.580000 ;
        RECT 1.030000 51.100000 2.230000 51.580000 ;
        RECT 1.030000 56.540000 2.230000 57.020000 ;
        RECT 4.895000 56.540000 6.260000 57.020000 ;
        RECT 1.030000 61.980000 2.230000 62.460000 ;
        RECT 4.895000 61.980000 6.260000 62.460000 ;
        RECT 1.030000 67.420000 2.230000 67.900000 ;
        RECT 4.895000 67.420000 6.260000 67.900000 ;
        RECT 1.030000 72.860000 2.230000 73.340000 ;
        RECT 4.895000 72.860000 6.260000 73.340000 ;
        RECT 4.895000 83.740000 6.260000 84.220000 ;
        RECT 1.030000 83.740000 2.230000 84.220000 ;
        RECT 4.895000 78.300000 6.260000 78.780000 ;
        RECT 1.030000 78.300000 2.230000 78.780000 ;
        RECT 1.030000 89.180000 2.230000 89.660000 ;
        RECT 4.895000 89.180000 6.260000 89.660000 ;
        RECT 1.030000 94.620000 2.230000 95.100000 ;
        RECT 4.895000 94.620000 6.260000 95.100000 ;
        RECT 37.790000 7.580000 38.990000 8.060000 ;
        RECT 37.790000 23.900000 38.990000 24.380000 ;
        RECT 37.790000 18.460000 38.990000 18.940000 ;
        RECT 37.790000 13.020000 38.990000 13.500000 ;
        RECT 37.790000 34.780000 38.990000 35.260000 ;
        RECT 37.790000 29.340000 38.990000 29.820000 ;
        RECT 37.790000 45.660000 38.990000 46.140000 ;
        RECT 37.790000 40.220000 38.990000 40.700000 ;
        RECT 37.790000 61.980000 38.990000 62.460000 ;
        RECT 37.790000 56.540000 38.990000 57.020000 ;
        RECT 37.790000 51.100000 38.990000 51.580000 ;
        RECT 37.790000 72.860000 38.990000 73.340000 ;
        RECT 37.790000 67.420000 38.990000 67.900000 ;
        RECT 37.790000 83.740000 38.990000 84.220000 ;
        RECT 37.790000 78.300000 38.990000 78.780000 ;
        RECT 37.790000 94.620000 38.990000 95.100000 ;
        RECT 37.790000 89.180000 38.990000 89.660000 ;
        RECT 1.030000 105.500000 2.230000 105.980000 ;
        RECT 4.895000 105.500000 6.260000 105.980000 ;
        RECT 1.030000 110.940000 2.230000 111.420000 ;
        RECT 4.895000 110.940000 6.260000 111.420000 ;
        RECT 4.895000 121.820000 6.260000 122.300000 ;
        RECT 1.030000 121.820000 2.230000 122.300000 ;
        RECT 4.895000 116.380000 6.260000 116.860000 ;
        RECT 1.030000 116.380000 2.230000 116.860000 ;
        RECT 1.030000 127.260000 2.230000 127.740000 ;
        RECT 4.895000 127.260000 6.260000 127.740000 ;
        RECT 1.030000 132.700000 2.230000 133.180000 ;
        RECT 4.895000 132.700000 6.260000 133.180000 ;
        RECT 4.895000 143.580000 6.260000 144.060000 ;
        RECT 1.030000 143.580000 2.230000 144.060000 ;
        RECT 4.895000 138.140000 6.260000 138.620000 ;
        RECT 1.030000 138.140000 2.230000 138.620000 ;
        RECT 1.030000 149.020000 2.230000 149.500000 ;
        RECT 4.895000 149.020000 6.260000 149.500000 ;
        RECT 1.030000 154.460000 2.230000 154.940000 ;
        RECT 4.895000 154.460000 6.260000 154.940000 ;
        RECT 1.030000 159.900000 2.230000 160.380000 ;
        RECT 4.895000 159.900000 6.260000 160.380000 ;
        RECT 1.030000 165.340000 2.230000 165.820000 ;
        RECT 4.895000 165.340000 6.260000 165.820000 ;
        RECT 1.030000 170.780000 2.230000 171.260000 ;
        RECT 4.895000 170.780000 6.260000 171.260000 ;
        RECT 4.895000 176.220000 6.260000 176.700000 ;
        RECT 1.030000 176.220000 2.230000 176.700000 ;
        RECT 1.030000 181.660000 2.230000 182.140000 ;
        RECT 4.895000 181.660000 6.260000 182.140000 ;
        RECT 1.030000 187.100000 2.230000 187.580000 ;
        RECT 4.895000 187.100000 6.260000 187.580000 ;
        RECT 4.895000 192.540000 6.260000 193.020000 ;
        RECT 1.030000 192.540000 2.230000 193.020000 ;
        RECT 37.790000 110.940000 38.990000 111.420000 ;
        RECT 37.790000 105.500000 38.990000 105.980000 ;
        RECT 37.790000 121.820000 38.990000 122.300000 ;
        RECT 37.790000 116.380000 38.990000 116.860000 ;
        RECT 37.790000 132.700000 38.990000 133.180000 ;
        RECT 37.790000 127.260000 38.990000 127.740000 ;
        RECT 37.790000 149.020000 38.990000 149.500000 ;
        RECT 37.790000 143.580000 38.990000 144.060000 ;
        RECT 37.790000 138.140000 38.990000 138.620000 ;
        RECT 37.790000 159.900000 38.990000 160.380000 ;
        RECT 37.790000 154.460000 38.990000 154.940000 ;
        RECT 37.790000 170.780000 38.990000 171.260000 ;
        RECT 37.790000 165.340000 38.990000 165.820000 ;
        RECT 37.790000 176.220000 38.990000 176.700000 ;
        RECT 37.790000 181.660000 38.990000 182.140000 ;
        RECT 37.790000 187.100000 38.990000 187.580000 ;
        RECT 37.790000 192.540000 38.990000 193.020000 ;
      LAYER met4 ;
        RECT 5.060000 1.050000 6.260000 198.020000 ;
        RECT 37.790000 0.000000 38.990000 200.260000 ;
        RECT 1.030000 0.000000 2.230000 200.260000 ;
        RECT 4.895000 100.060000 6.260000 100.540000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
        RECT 4.895000 29.340000 6.260000 29.820000 ;
        RECT 4.895000 34.780000 6.260000 35.260000 ;
        RECT 4.895000 40.220000 6.260000 40.700000 ;
        RECT 4.895000 45.660000 6.260000 46.140000 ;
        RECT 4.895000 51.100000 6.260000 51.580000 ;
        RECT 4.895000 56.540000 6.260000 57.020000 ;
        RECT 4.895000 61.980000 6.260000 62.460000 ;
        RECT 4.895000 67.420000 6.260000 67.900000 ;
        RECT 4.895000 72.860000 6.260000 73.340000 ;
        RECT 4.895000 83.740000 6.260000 84.220000 ;
        RECT 4.895000 78.300000 6.260000 78.780000 ;
        RECT 4.895000 89.180000 6.260000 89.660000 ;
        RECT 4.895000 94.620000 6.260000 95.100000 ;
        RECT 4.895000 105.500000 6.260000 105.980000 ;
        RECT 4.895000 110.940000 6.260000 111.420000 ;
        RECT 4.895000 121.820000 6.260000 122.300000 ;
        RECT 4.895000 116.380000 6.260000 116.860000 ;
        RECT 4.895000 127.260000 6.260000 127.740000 ;
        RECT 4.895000 132.700000 6.260000 133.180000 ;
        RECT 4.895000 143.580000 6.260000 144.060000 ;
        RECT 4.895000 138.140000 6.260000 138.620000 ;
        RECT 4.895000 149.020000 6.260000 149.500000 ;
        RECT 4.895000 154.460000 6.260000 154.940000 ;
        RECT 4.895000 159.900000 6.260000 160.380000 ;
        RECT 4.895000 165.340000 6.260000 165.820000 ;
        RECT 4.895000 170.780000 6.260000 171.260000 ;
        RECT 4.895000 176.220000 6.260000 176.700000 ;
        RECT 4.895000 181.660000 6.260000 182.140000 ;
        RECT 4.895000 187.100000 6.260000 187.580000 ;
        RECT 4.895000 192.540000 6.260000 193.020000 ;
    END
# end of P/G power stripe data as pin

  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 40.020000 200.260000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 40.020000 200.260000 ;
    LAYER met2 ;
      RECT 35.060000 199.420000 40.020000 200.260000 ;
      RECT 33.220000 199.420000 34.400000 200.260000 ;
      RECT 31.840000 199.420000 32.560000 200.260000 ;
      RECT 30.460000 199.420000 31.180000 200.260000 ;
      RECT 29.080000 199.420000 29.800000 200.260000 ;
      RECT 27.700000 199.420000 28.420000 200.260000 ;
      RECT 25.860000 199.420000 27.040000 200.260000 ;
      RECT 24.480000 199.420000 25.200000 200.260000 ;
      RECT 23.100000 199.420000 23.820000 200.260000 ;
      RECT 21.720000 199.420000 22.440000 200.260000 ;
      RECT 19.880000 199.420000 21.060000 200.260000 ;
      RECT 18.500000 199.420000 19.220000 200.260000 ;
      RECT 17.120000 199.420000 17.840000 200.260000 ;
      RECT 15.740000 199.420000 16.460000 200.260000 ;
      RECT 14.360000 199.420000 15.080000 200.260000 ;
      RECT 12.980000 199.420000 13.700000 200.260000 ;
      RECT 11.140000 199.420000 12.320000 200.260000 ;
      RECT 9.760000 199.420000 10.480000 200.260000 ;
      RECT 8.380000 199.420000 9.100000 200.260000 ;
      RECT 7.000000 199.420000 7.720000 200.260000 ;
      RECT 5.620000 199.420000 6.340000 200.260000 ;
      RECT 0.000000 199.420000 4.960000 200.260000 ;
      RECT 0.000000 0.840000 40.020000 199.420000 ;
      RECT 35.060000 0.000000 40.020000 0.840000 ;
      RECT 33.220000 0.000000 34.400000 0.840000 ;
      RECT 31.840000 0.000000 32.560000 0.840000 ;
      RECT 30.460000 0.000000 31.180000 0.840000 ;
      RECT 29.080000 0.000000 29.800000 0.840000 ;
      RECT 27.700000 0.000000 28.420000 0.840000 ;
      RECT 25.860000 0.000000 27.040000 0.840000 ;
      RECT 24.480000 0.000000 25.200000 0.840000 ;
      RECT 23.100000 0.000000 23.820000 0.840000 ;
      RECT 21.720000 0.000000 22.440000 0.840000 ;
      RECT 19.880000 0.000000 21.060000 0.840000 ;
      RECT 18.500000 0.000000 19.220000 0.840000 ;
      RECT 17.120000 0.000000 17.840000 0.840000 ;
      RECT 15.740000 0.000000 16.460000 0.840000 ;
      RECT 14.360000 0.000000 15.080000 0.840000 ;
      RECT 12.980000 0.000000 13.700000 0.840000 ;
      RECT 11.140000 0.000000 12.320000 0.840000 ;
      RECT 9.760000 0.000000 10.480000 0.840000 ;
      RECT 8.380000 0.000000 9.100000 0.840000 ;
      RECT 7.000000 0.000000 7.720000 0.840000 ;
      RECT 5.620000 0.000000 6.340000 0.840000 ;
      RECT 0.000000 0.000000 4.960000 0.840000 ;
    LAYER met3 ;
      RECT 0.000000 198.320000 40.020000 200.260000 ;
      RECT 1.000000 194.250000 40.020000 194.720000 ;
      RECT 1.000000 193.880000 39.020000 194.250000 ;
      RECT 0.000000 193.320000 39.020000 193.880000 ;
      RECT 0.000000 193.030000 0.730000 193.320000 ;
      RECT 39.290000 192.240000 40.020000 193.270000 ;
      RECT 6.560000 192.240000 37.490000 193.320000 ;
      RECT 2.530000 192.240000 4.595000 193.320000 ;
      RECT 1.000000 192.050000 40.020000 192.240000 ;
      RECT 0.000000 191.810000 40.020000 192.050000 ;
      RECT 1.000000 190.830000 40.020000 191.810000 ;
      RECT 0.000000 190.600000 40.020000 190.830000 ;
      RECT 37.490000 190.590000 40.020000 190.600000 ;
      RECT 0.000000 189.980000 2.530000 190.600000 ;
      RECT 37.490000 189.610000 39.020000 190.590000 ;
      RECT 37.490000 189.520000 40.020000 189.610000 ;
      RECT 8.560000 189.520000 35.690000 190.600000 ;
      RECT 4.330000 189.520000 6.760000 190.600000 ;
      RECT 1.000000 189.520000 2.530000 189.980000 ;
      RECT 1.000000 189.000000 40.020000 189.520000 ;
      RECT 0.000000 188.760000 40.020000 189.000000 ;
      RECT 1.000000 187.880000 40.020000 188.760000 ;
      RECT 39.290000 186.930000 40.020000 187.880000 ;
      RECT 0.000000 186.930000 0.730000 187.780000 ;
      RECT 6.560000 186.800000 37.490000 187.880000 ;
      RECT 2.530000 186.800000 4.595000 187.880000 ;
      RECT 1.000000 185.950000 39.020000 186.800000 ;
      RECT 0.000000 185.710000 40.020000 185.950000 ;
      RECT 1.000000 185.160000 40.020000 185.710000 ;
      RECT 1.000000 184.730000 2.530000 185.160000 ;
      RECT 37.490000 184.080000 40.020000 185.160000 ;
      RECT 8.560000 184.080000 35.690000 185.160000 ;
      RECT 4.330000 184.080000 6.760000 185.160000 ;
      RECT 0.000000 184.080000 2.530000 184.730000 ;
      RECT 0.000000 183.880000 40.020000 184.080000 ;
      RECT 1.000000 183.270000 40.020000 183.880000 ;
      RECT 1.000000 182.900000 39.020000 183.270000 ;
      RECT 0.000000 182.660000 39.020000 182.900000 ;
      RECT 1.000000 182.440000 39.020000 182.660000 ;
      RECT 0.000000 181.440000 0.730000 181.680000 ;
      RECT 39.290000 181.360000 40.020000 182.290000 ;
      RECT 6.560000 181.360000 37.490000 182.440000 ;
      RECT 2.530000 181.360000 4.595000 182.440000 ;
      RECT 1.000000 180.460000 40.020000 181.360000 ;
      RECT 0.000000 179.720000 40.020000 180.460000 ;
      RECT 37.490000 179.610000 40.020000 179.720000 ;
      RECT 0.000000 179.610000 2.530000 179.720000 ;
      RECT 37.490000 178.640000 39.020000 179.610000 ;
      RECT 8.560000 178.640000 35.690000 179.720000 ;
      RECT 4.330000 178.640000 6.760000 179.720000 ;
      RECT 1.000000 178.640000 2.530000 179.610000 ;
      RECT 1.000000 178.630000 39.020000 178.640000 ;
      RECT 0.000000 178.390000 40.020000 178.630000 ;
      RECT 1.000000 177.410000 40.020000 178.390000 ;
      RECT 0.000000 177.000000 40.020000 177.410000 ;
      RECT 0.000000 176.560000 0.730000 177.000000 ;
      RECT 39.290000 175.950000 40.020000 177.000000 ;
      RECT 6.560000 175.920000 37.490000 177.000000 ;
      RECT 2.530000 175.920000 4.595000 177.000000 ;
      RECT 1.000000 175.580000 39.020000 175.920000 ;
      RECT 0.000000 175.340000 39.020000 175.580000 ;
      RECT 1.000000 174.970000 39.020000 175.340000 ;
      RECT 1.000000 174.360000 40.020000 174.970000 ;
      RECT 0.000000 174.280000 40.020000 174.360000 ;
      RECT 0.000000 173.510000 2.530000 174.280000 ;
      RECT 37.490000 173.200000 40.020000 174.280000 ;
      RECT 8.560000 173.200000 35.690000 174.280000 ;
      RECT 4.330000 173.200000 6.760000 174.280000 ;
      RECT 1.000000 173.200000 2.530000 173.510000 ;
      RECT 1.000000 172.530000 40.020000 173.200000 ;
      RECT 0.000000 172.290000 40.020000 172.530000 ;
      RECT 1.000000 171.560000 39.020000 172.290000 ;
      RECT 39.290000 170.480000 40.020000 171.310000 ;
      RECT 6.560000 170.480000 37.490000 171.560000 ;
      RECT 2.530000 170.480000 4.595000 171.560000 ;
      RECT 0.000000 170.480000 0.730000 171.310000 ;
      RECT 0.000000 170.460000 40.020000 170.480000 ;
      RECT 1.000000 169.480000 40.020000 170.460000 ;
      RECT 0.000000 169.240000 40.020000 169.480000 ;
      RECT 1.000000 168.840000 40.020000 169.240000 ;
      RECT 37.490000 168.630000 40.020000 168.840000 ;
      RECT 1.000000 168.260000 2.530000 168.840000 ;
      RECT 0.000000 168.020000 2.530000 168.260000 ;
      RECT 37.490000 167.760000 39.020000 168.630000 ;
      RECT 8.560000 167.760000 35.690000 168.840000 ;
      RECT 4.330000 167.760000 6.760000 168.840000 ;
      RECT 1.000000 167.760000 2.530000 168.020000 ;
      RECT 1.000000 167.650000 39.020000 167.760000 ;
      RECT 1.000000 167.040000 40.020000 167.650000 ;
      RECT 0.000000 166.190000 40.020000 167.040000 ;
      RECT 1.000000 166.120000 40.020000 166.190000 ;
      RECT 39.290000 165.040000 40.020000 166.120000 ;
      RECT 6.560000 165.040000 37.490000 166.120000 ;
      RECT 2.530000 165.040000 4.595000 166.120000 ;
      RECT 0.000000 165.040000 0.730000 165.210000 ;
      RECT 0.000000 164.970000 40.020000 165.040000 ;
      RECT 1.000000 163.990000 39.020000 164.970000 ;
      RECT 0.000000 163.400000 40.020000 163.990000 ;
      RECT 0.000000 163.140000 2.530000 163.400000 ;
      RECT 37.490000 162.320000 40.020000 163.400000 ;
      RECT 8.560000 162.320000 35.690000 163.400000 ;
      RECT 4.330000 162.320000 6.760000 163.400000 ;
      RECT 1.000000 162.320000 2.530000 163.140000 ;
      RECT 1.000000 162.160000 40.020000 162.320000 ;
      RECT 0.000000 161.920000 40.020000 162.160000 ;
      RECT 1.000000 161.310000 40.020000 161.920000 ;
      RECT 1.000000 160.940000 39.020000 161.310000 ;
      RECT 0.000000 160.680000 39.020000 160.940000 ;
      RECT 0.000000 160.090000 0.730000 160.680000 ;
      RECT 39.290000 159.600000 40.020000 160.330000 ;
      RECT 6.560000 159.600000 37.490000 160.680000 ;
      RECT 2.530000 159.600000 4.595000 160.680000 ;
      RECT 1.000000 159.110000 40.020000 159.600000 ;
      RECT 0.000000 158.870000 40.020000 159.110000 ;
      RECT 1.000000 157.960000 40.020000 158.870000 ;
      RECT 1.000000 157.890000 2.530000 157.960000 ;
      RECT 37.490000 157.650000 40.020000 157.960000 ;
      RECT 0.000000 157.040000 2.530000 157.890000 ;
      RECT 37.490000 156.880000 39.020000 157.650000 ;
      RECT 8.560000 156.880000 35.690000 157.960000 ;
      RECT 4.330000 156.880000 6.760000 157.960000 ;
      RECT 1.000000 156.880000 2.530000 157.040000 ;
      RECT 1.000000 156.670000 39.020000 156.880000 ;
      RECT 1.000000 156.060000 40.020000 156.670000 ;
      RECT 0.000000 155.820000 40.020000 156.060000 ;
      RECT 1.000000 155.240000 40.020000 155.820000 ;
      RECT 0.000000 154.600000 0.730000 154.840000 ;
      RECT 39.290000 154.160000 40.020000 155.240000 ;
      RECT 6.560000 154.160000 37.490000 155.240000 ;
      RECT 2.530000 154.160000 4.595000 155.240000 ;
      RECT 1.000000 153.990000 40.020000 154.160000 ;
      RECT 1.000000 153.620000 39.020000 153.990000 ;
      RECT 0.000000 153.010000 39.020000 153.620000 ;
      RECT 0.000000 152.770000 40.020000 153.010000 ;
      RECT 1.000000 152.520000 40.020000 152.770000 ;
      RECT 1.000000 151.790000 2.530000 152.520000 ;
      RECT 0.000000 151.550000 2.530000 151.790000 ;
      RECT 37.490000 151.440000 40.020000 152.520000 ;
      RECT 8.560000 151.440000 35.690000 152.520000 ;
      RECT 4.330000 151.440000 6.760000 152.520000 ;
      RECT 1.000000 151.440000 2.530000 151.550000 ;
      RECT 1.000000 150.570000 40.020000 151.440000 ;
      RECT 0.000000 150.330000 40.020000 150.570000 ;
      RECT 0.000000 149.800000 39.020000 150.330000 ;
      RECT 0.000000 149.720000 0.730000 149.800000 ;
      RECT 39.290000 148.720000 40.020000 149.350000 ;
      RECT 6.560000 148.720000 37.490000 149.800000 ;
      RECT 2.530000 148.720000 4.595000 149.800000 ;
      RECT 0.000000 148.720000 0.730000 148.740000 ;
      RECT 0.000000 148.500000 40.020000 148.720000 ;
      RECT 1.000000 147.520000 40.020000 148.500000 ;
      RECT 0.000000 147.080000 40.020000 147.520000 ;
      RECT 0.000000 146.670000 2.530000 147.080000 ;
      RECT 37.490000 146.060000 40.020000 147.080000 ;
      RECT 37.490000 146.000000 39.020000 146.060000 ;
      RECT 8.560000 146.000000 35.690000 147.080000 ;
      RECT 4.330000 146.000000 6.760000 147.080000 ;
      RECT 1.000000 146.000000 2.530000 146.670000 ;
      RECT 1.000000 145.690000 39.020000 146.000000 ;
      RECT 0.000000 145.450000 39.020000 145.690000 ;
      RECT 1.000000 145.080000 39.020000 145.450000 ;
      RECT 1.000000 144.470000 40.020000 145.080000 ;
      RECT 0.000000 144.360000 40.020000 144.470000 ;
      RECT 0.000000 144.230000 0.730000 144.360000 ;
      RECT 39.290000 143.280000 40.020000 144.360000 ;
      RECT 6.560000 143.280000 37.490000 144.360000 ;
      RECT 2.530000 143.280000 4.595000 144.360000 ;
      RECT 1.000000 143.250000 40.020000 143.280000 ;
      RECT 0.000000 142.400000 40.020000 143.250000 ;
      RECT 1.000000 141.640000 39.020000 142.400000 ;
      RECT 37.490000 141.420000 39.020000 141.640000 ;
      RECT 1.000000 141.420000 2.530000 141.640000 ;
      RECT 0.000000 141.180000 2.530000 141.420000 ;
      RECT 37.490000 140.560000 40.020000 141.420000 ;
      RECT 8.560000 140.560000 35.690000 141.640000 ;
      RECT 4.330000 140.560000 6.760000 141.640000 ;
      RECT 1.000000 140.560000 2.530000 141.180000 ;
      RECT 1.000000 140.200000 40.020000 140.560000 ;
      RECT 0.000000 139.350000 40.020000 140.200000 ;
      RECT 1.000000 138.920000 40.020000 139.350000 ;
      RECT 39.290000 138.740000 40.020000 138.920000 ;
      RECT 0.000000 138.130000 0.730000 138.370000 ;
      RECT 6.560000 137.840000 37.490000 138.920000 ;
      RECT 2.530000 137.840000 4.595000 138.920000 ;
      RECT 1.000000 137.760000 39.020000 137.840000 ;
      RECT 1.000000 137.150000 40.020000 137.760000 ;
      RECT 0.000000 136.300000 40.020000 137.150000 ;
      RECT 1.000000 136.200000 40.020000 136.300000 ;
      RECT 1.000000 135.320000 2.530000 136.200000 ;
      RECT 37.490000 135.120000 40.020000 136.200000 ;
      RECT 8.560000 135.120000 35.690000 136.200000 ;
      RECT 4.330000 135.120000 6.760000 136.200000 ;
      RECT 0.000000 135.120000 2.530000 135.320000 ;
      RECT 0.000000 135.080000 40.020000 135.120000 ;
      RECT 1.000000 134.100000 39.020000 135.080000 ;
      RECT 0.000000 133.480000 40.020000 134.100000 ;
      RECT 0.000000 133.250000 0.730000 133.480000 ;
      RECT 39.290000 132.400000 40.020000 133.480000 ;
      RECT 6.560000 132.400000 37.490000 133.480000 ;
      RECT 2.530000 132.400000 4.595000 133.480000 ;
      RECT 1.000000 132.270000 40.020000 132.400000 ;
      RECT 0.000000 132.030000 40.020000 132.270000 ;
      RECT 1.000000 131.420000 40.020000 132.030000 ;
      RECT 1.000000 131.050000 39.020000 131.420000 ;
      RECT 0.000000 130.810000 39.020000 131.050000 ;
      RECT 1.000000 130.760000 39.020000 130.810000 ;
      RECT 37.490000 130.440000 39.020000 130.760000 ;
      RECT 1.000000 129.830000 2.530000 130.760000 ;
      RECT 37.490000 129.680000 40.020000 130.440000 ;
      RECT 8.560000 129.680000 35.690000 130.760000 ;
      RECT 4.330000 129.680000 6.760000 130.760000 ;
      RECT 0.000000 129.680000 2.530000 129.830000 ;
      RECT 0.000000 128.980000 40.020000 129.680000 ;
      RECT 1.000000 128.040000 40.020000 128.980000 ;
      RECT 39.290000 127.760000 40.020000 128.040000 ;
      RECT 0.000000 127.760000 0.730000 128.000000 ;
      RECT 6.560000 126.960000 37.490000 128.040000 ;
      RECT 2.530000 126.960000 4.595000 128.040000 ;
      RECT 1.000000 126.780000 39.020000 126.960000 ;
      RECT 0.000000 125.930000 40.020000 126.780000 ;
      RECT 1.000000 125.320000 40.020000 125.930000 ;
      RECT 1.000000 124.950000 2.530000 125.320000 ;
      RECT 0.000000 124.710000 2.530000 124.950000 ;
      RECT 37.490000 124.240000 40.020000 125.320000 ;
      RECT 8.560000 124.240000 35.690000 125.320000 ;
      RECT 4.330000 124.240000 6.760000 125.320000 ;
      RECT 1.000000 124.240000 2.530000 124.710000 ;
      RECT 1.000000 124.100000 40.020000 124.240000 ;
      RECT 1.000000 123.730000 39.020000 124.100000 ;
      RECT 0.000000 123.120000 39.020000 123.730000 ;
      RECT 0.000000 122.880000 40.020000 123.120000 ;
      RECT 1.000000 122.600000 40.020000 122.880000 ;
      RECT 0.000000 121.660000 0.730000 121.900000 ;
      RECT 39.290000 121.520000 40.020000 122.600000 ;
      RECT 6.560000 121.520000 37.490000 122.600000 ;
      RECT 2.530000 121.520000 4.595000 122.600000 ;
      RECT 1.000000 120.680000 40.020000 121.520000 ;
      RECT 0.000000 120.440000 40.020000 120.680000 ;
      RECT 0.000000 119.880000 39.020000 120.440000 ;
      RECT 0.000000 119.830000 2.530000 119.880000 ;
      RECT 37.490000 119.460000 39.020000 119.880000 ;
      RECT 1.000000 118.850000 2.530000 119.830000 ;
      RECT 37.490000 118.800000 40.020000 119.460000 ;
      RECT 8.560000 118.800000 35.690000 119.880000 ;
      RECT 4.330000 118.800000 6.760000 119.880000 ;
      RECT 0.000000 118.800000 2.530000 118.850000 ;
      RECT 0.000000 118.610000 40.020000 118.800000 ;
      RECT 1.000000 117.630000 40.020000 118.610000 ;
      RECT 0.000000 117.390000 40.020000 117.630000 ;
      RECT 1.000000 117.160000 40.020000 117.390000 ;
      RECT 39.290000 116.780000 40.020000 117.160000 ;
      RECT 6.560000 116.080000 37.490000 117.160000 ;
      RECT 2.530000 116.080000 4.595000 117.160000 ;
      RECT 0.000000 116.080000 0.730000 116.410000 ;
      RECT 0.000000 115.800000 39.020000 116.080000 ;
      RECT 0.000000 115.560000 40.020000 115.800000 ;
      RECT 1.000000 114.580000 40.020000 115.560000 ;
      RECT 0.000000 114.440000 40.020000 114.580000 ;
      RECT 0.000000 114.340000 2.530000 114.440000 ;
      RECT 37.490000 113.360000 40.020000 114.440000 ;
      RECT 8.560000 113.360000 35.690000 114.440000 ;
      RECT 4.330000 113.360000 6.760000 114.440000 ;
      RECT 1.000000 113.360000 2.530000 114.340000 ;
      RECT 0.000000 113.120000 40.020000 113.360000 ;
      RECT 0.000000 112.510000 39.020000 113.120000 ;
      RECT 1.000000 112.140000 39.020000 112.510000 ;
      RECT 1.000000 111.720000 40.020000 112.140000 ;
      RECT 0.000000 111.290000 0.730000 111.530000 ;
      RECT 39.290000 110.640000 40.020000 111.720000 ;
      RECT 6.560000 110.640000 37.490000 111.720000 ;
      RECT 2.530000 110.640000 4.595000 111.720000 ;
      RECT 1.000000 110.310000 40.020000 110.640000 ;
      RECT 0.000000 109.460000 40.020000 110.310000 ;
      RECT 1.000000 109.000000 39.020000 109.460000 ;
      RECT 37.490000 108.480000 39.020000 109.000000 ;
      RECT 1.000000 108.480000 2.530000 109.000000 ;
      RECT 0.000000 108.240000 2.530000 108.480000 ;
      RECT 37.490000 107.920000 40.020000 108.480000 ;
      RECT 8.560000 107.920000 35.690000 109.000000 ;
      RECT 4.330000 107.920000 6.760000 109.000000 ;
      RECT 1.000000 107.920000 2.530000 108.240000 ;
      RECT 1.000000 107.260000 40.020000 107.920000 ;
      RECT 0.000000 106.410000 40.020000 107.260000 ;
      RECT 1.000000 106.280000 40.020000 106.410000 ;
      RECT 39.290000 105.800000 40.020000 106.280000 ;
      RECT 6.560000 105.200000 37.490000 106.280000 ;
      RECT 2.530000 105.200000 4.595000 106.280000 ;
      RECT 0.000000 105.200000 0.730000 105.430000 ;
      RECT 0.000000 105.190000 39.020000 105.200000 ;
      RECT 1.000000 104.820000 39.020000 105.190000 ;
      RECT 1.000000 104.210000 40.020000 104.820000 ;
      RECT 0.000000 103.970000 40.020000 104.210000 ;
      RECT 1.000000 103.560000 40.020000 103.970000 ;
      RECT 1.000000 102.990000 2.530000 103.560000 ;
      RECT 37.490000 102.480000 40.020000 103.560000 ;
      RECT 8.560000 102.480000 35.690000 103.560000 ;
      RECT 4.330000 102.480000 6.760000 103.560000 ;
      RECT 0.000000 102.480000 2.530000 102.990000 ;
      RECT 0.000000 102.140000 40.020000 102.480000 ;
      RECT 1.000000 101.160000 39.020000 102.140000 ;
      RECT 0.000000 100.920000 40.020000 101.160000 ;
      RECT 1.000000 100.840000 40.020000 100.920000 ;
      RECT 39.290000 99.760000 40.020000 100.840000 ;
      RECT 6.560000 99.760000 37.490000 100.840000 ;
      RECT 2.530000 99.760000 4.595000 100.840000 ;
      RECT 0.000000 99.760000 0.730000 99.940000 ;
      RECT 0.000000 99.090000 40.020000 99.760000 ;
      RECT 1.000000 98.120000 40.020000 99.090000 ;
      RECT 1.000000 98.110000 2.530000 98.120000 ;
      RECT 37.490000 97.870000 40.020000 98.120000 ;
      RECT 0.000000 97.870000 2.530000 98.110000 ;
      RECT 37.490000 97.040000 39.020000 97.870000 ;
      RECT 8.560000 97.040000 35.690000 98.120000 ;
      RECT 4.330000 97.040000 6.760000 98.120000 ;
      RECT 1.000000 97.040000 2.530000 97.870000 ;
      RECT 1.000000 96.890000 39.020000 97.040000 ;
      RECT 0.000000 96.040000 40.020000 96.890000 ;
      RECT 1.000000 95.400000 40.020000 96.040000 ;
      RECT 0.000000 94.820000 0.730000 95.060000 ;
      RECT 39.290000 94.320000 40.020000 95.400000 ;
      RECT 6.560000 94.320000 37.490000 95.400000 ;
      RECT 2.530000 94.320000 4.595000 95.400000 ;
      RECT 1.000000 94.210000 40.020000 94.320000 ;
      RECT 1.000000 93.840000 39.020000 94.210000 ;
      RECT 0.000000 93.600000 39.020000 93.840000 ;
      RECT 1.000000 93.230000 39.020000 93.600000 ;
      RECT 1.000000 92.680000 40.020000 93.230000 ;
      RECT 1.000000 92.620000 2.530000 92.680000 ;
      RECT 0.000000 91.770000 2.530000 92.620000 ;
      RECT 37.490000 91.600000 40.020000 92.680000 ;
      RECT 8.560000 91.600000 35.690000 92.680000 ;
      RECT 4.330000 91.600000 6.760000 92.680000 ;
      RECT 1.000000 91.600000 2.530000 91.770000 ;
      RECT 1.000000 90.790000 40.020000 91.600000 ;
      RECT 0.000000 90.550000 40.020000 90.790000 ;
      RECT 1.000000 89.960000 39.020000 90.550000 ;
      RECT 39.290000 88.880000 40.020000 89.570000 ;
      RECT 6.560000 88.880000 37.490000 89.960000 ;
      RECT 2.530000 88.880000 4.595000 89.960000 ;
      RECT 0.000000 88.880000 0.730000 89.570000 ;
      RECT 0.000000 88.720000 40.020000 88.880000 ;
      RECT 1.000000 87.740000 40.020000 88.720000 ;
      RECT 0.000000 87.500000 40.020000 87.740000 ;
      RECT 1.000000 87.240000 40.020000 87.500000 ;
      RECT 37.490000 86.890000 40.020000 87.240000 ;
      RECT 1.000000 86.520000 2.530000 87.240000 ;
      RECT 37.490000 86.160000 39.020000 86.890000 ;
      RECT 8.560000 86.160000 35.690000 87.240000 ;
      RECT 4.330000 86.160000 6.760000 87.240000 ;
      RECT 0.000000 86.160000 2.530000 86.520000 ;
      RECT 0.000000 85.910000 39.020000 86.160000 ;
      RECT 0.000000 85.670000 40.020000 85.910000 ;
      RECT 1.000000 84.690000 40.020000 85.670000 ;
      RECT 0.000000 84.520000 40.020000 84.690000 ;
      RECT 0.000000 84.450000 0.730000 84.520000 ;
      RECT 39.290000 83.440000 40.020000 84.520000 ;
      RECT 6.560000 83.440000 37.490000 84.520000 ;
      RECT 2.530000 83.440000 4.595000 84.520000 ;
      RECT 0.000000 83.440000 0.730000 83.470000 ;
      RECT 0.000000 83.230000 40.020000 83.440000 ;
      RECT 0.000000 82.620000 39.020000 83.230000 ;
      RECT 1.000000 82.250000 39.020000 82.620000 ;
      RECT 1.000000 81.800000 40.020000 82.250000 ;
      RECT 1.000000 81.640000 2.530000 81.800000 ;
      RECT 0.000000 81.400000 2.530000 81.640000 ;
      RECT 37.490000 80.720000 40.020000 81.800000 ;
      RECT 8.560000 80.720000 35.690000 81.800000 ;
      RECT 4.330000 80.720000 6.760000 81.800000 ;
      RECT 1.000000 80.720000 2.530000 81.400000 ;
      RECT 1.000000 80.420000 40.020000 80.720000 ;
      RECT 0.000000 80.180000 40.020000 80.420000 ;
      RECT 1.000000 79.570000 40.020000 80.180000 ;
      RECT 1.000000 79.200000 39.020000 79.570000 ;
      RECT 0.000000 79.080000 39.020000 79.200000 ;
      RECT 0.000000 78.350000 0.730000 79.080000 ;
      RECT 39.290000 78.000000 40.020000 78.590000 ;
      RECT 6.560000 78.000000 37.490000 79.080000 ;
      RECT 2.530000 78.000000 4.595000 79.080000 ;
      RECT 1.000000 77.370000 40.020000 78.000000 ;
      RECT 0.000000 77.130000 40.020000 77.370000 ;
      RECT 1.000000 76.360000 40.020000 77.130000 ;
      RECT 1.000000 76.150000 2.530000 76.360000 ;
      RECT 37.490000 75.910000 40.020000 76.360000 ;
      RECT 0.000000 75.300000 2.530000 76.150000 ;
      RECT 37.490000 75.280000 39.020000 75.910000 ;
      RECT 8.560000 75.280000 35.690000 76.360000 ;
      RECT 4.330000 75.280000 6.760000 76.360000 ;
      RECT 1.000000 75.280000 2.530000 75.300000 ;
      RECT 1.000000 74.930000 39.020000 75.280000 ;
      RECT 1.000000 74.320000 40.020000 74.930000 ;
      RECT 0.000000 74.080000 40.020000 74.320000 ;
      RECT 1.000000 73.640000 40.020000 74.080000 ;
      RECT 39.290000 72.560000 40.020000 73.640000 ;
      RECT 6.560000 72.560000 37.490000 73.640000 ;
      RECT 2.530000 72.560000 4.595000 73.640000 ;
      RECT 0.000000 72.560000 0.730000 73.100000 ;
      RECT 0.000000 72.250000 40.020000 72.560000 ;
      RECT 1.000000 71.270000 39.020000 72.250000 ;
      RECT 0.000000 71.030000 40.020000 71.270000 ;
      RECT 1.000000 70.920000 40.020000 71.030000 ;
      RECT 1.000000 70.050000 2.530000 70.920000 ;
      RECT 37.490000 69.840000 40.020000 70.920000 ;
      RECT 8.560000 69.840000 35.690000 70.920000 ;
      RECT 4.330000 69.840000 6.760000 70.920000 ;
      RECT 0.000000 69.840000 2.530000 70.050000 ;
      RECT 0.000000 69.200000 40.020000 69.840000 ;
      RECT 1.000000 68.590000 40.020000 69.200000 ;
      RECT 1.000000 68.220000 39.020000 68.590000 ;
      RECT 0.000000 68.200000 39.020000 68.220000 ;
      RECT 0.000000 67.980000 0.730000 68.200000 ;
      RECT 39.290000 67.120000 40.020000 67.610000 ;
      RECT 6.560000 67.120000 37.490000 68.200000 ;
      RECT 2.530000 67.120000 4.595000 68.200000 ;
      RECT 1.000000 67.000000 40.020000 67.120000 ;
      RECT 0.000000 66.760000 40.020000 67.000000 ;
      RECT 1.000000 65.780000 40.020000 66.760000 ;
      RECT 0.000000 65.480000 40.020000 65.780000 ;
      RECT 37.490000 64.930000 40.020000 65.480000 ;
      RECT 0.000000 64.930000 2.530000 65.480000 ;
      RECT 37.490000 64.400000 39.020000 64.930000 ;
      RECT 8.560000 64.400000 35.690000 65.480000 ;
      RECT 4.330000 64.400000 6.760000 65.480000 ;
      RECT 1.000000 64.400000 2.530000 64.930000 ;
      RECT 1.000000 63.950000 39.020000 64.400000 ;
      RECT 0.000000 63.710000 40.020000 63.950000 ;
      RECT 1.000000 62.760000 40.020000 63.710000 ;
      RECT 0.000000 61.880000 0.730000 62.730000 ;
      RECT 39.290000 61.680000 40.020000 62.760000 ;
      RECT 6.560000 61.680000 37.490000 62.760000 ;
      RECT 2.530000 61.680000 4.595000 62.760000 ;
      RECT 1.000000 61.270000 40.020000 61.680000 ;
      RECT 1.000000 60.900000 39.020000 61.270000 ;
      RECT 0.000000 60.660000 39.020000 60.900000 ;
      RECT 1.000000 60.290000 39.020000 60.660000 ;
      RECT 1.000000 60.040000 40.020000 60.290000 ;
      RECT 1.000000 59.680000 2.530000 60.040000 ;
      RECT 37.490000 58.960000 40.020000 60.040000 ;
      RECT 8.560000 58.960000 35.690000 60.040000 ;
      RECT 4.330000 58.960000 6.760000 60.040000 ;
      RECT 0.000000 58.960000 2.530000 59.680000 ;
      RECT 0.000000 58.830000 40.020000 58.960000 ;
      RECT 1.000000 57.850000 40.020000 58.830000 ;
      RECT 0.000000 57.610000 40.020000 57.850000 ;
      RECT 1.000000 57.320000 39.020000 57.610000 ;
      RECT 39.290000 56.240000 40.020000 56.630000 ;
      RECT 6.560000 56.240000 37.490000 57.320000 ;
      RECT 2.530000 56.240000 4.595000 57.320000 ;
      RECT 0.000000 56.240000 0.730000 56.630000 ;
      RECT 0.000000 55.780000 40.020000 56.240000 ;
      RECT 1.000000 54.800000 40.020000 55.780000 ;
      RECT 0.000000 54.600000 40.020000 54.800000 ;
      RECT 0.000000 54.560000 2.530000 54.600000 ;
      RECT 37.490000 53.950000 40.020000 54.600000 ;
      RECT 1.000000 53.580000 2.530000 54.560000 ;
      RECT 37.490000 53.520000 39.020000 53.950000 ;
      RECT 8.560000 53.520000 35.690000 54.600000 ;
      RECT 4.330000 53.520000 6.760000 54.600000 ;
      RECT 0.000000 53.520000 2.530000 53.580000 ;
      RECT 0.000000 53.340000 39.020000 53.520000 ;
      RECT 1.000000 52.970000 39.020000 53.340000 ;
      RECT 1.000000 52.360000 40.020000 52.970000 ;
      RECT 0.000000 51.880000 40.020000 52.360000 ;
      RECT 0.000000 51.510000 0.730000 51.880000 ;
      RECT 39.290000 50.800000 40.020000 51.880000 ;
      RECT 6.560000 50.800000 37.490000 51.880000 ;
      RECT 2.530000 50.800000 4.595000 51.880000 ;
      RECT 1.000000 50.530000 40.020000 50.800000 ;
      RECT 0.000000 50.290000 40.020000 50.530000 ;
      RECT 1.000000 49.680000 40.020000 50.290000 ;
      RECT 1.000000 49.310000 39.020000 49.680000 ;
      RECT 0.000000 49.160000 39.020000 49.310000 ;
      RECT 37.490000 48.700000 39.020000 49.160000 ;
      RECT 0.000000 48.460000 2.530000 49.160000 ;
      RECT 37.490000 48.080000 40.020000 48.700000 ;
      RECT 8.560000 48.080000 35.690000 49.160000 ;
      RECT 4.330000 48.080000 6.760000 49.160000 ;
      RECT 1.000000 48.080000 2.530000 48.460000 ;
      RECT 1.000000 47.480000 40.020000 48.080000 ;
      RECT 0.000000 47.240000 40.020000 47.480000 ;
      RECT 1.000000 46.440000 40.020000 47.240000 ;
      RECT 39.290000 46.020000 40.020000 46.440000 ;
      RECT 0.000000 45.410000 0.730000 46.260000 ;
      RECT 6.560000 45.360000 37.490000 46.440000 ;
      RECT 2.530000 45.360000 4.595000 46.440000 ;
      RECT 1.000000 45.040000 39.020000 45.360000 ;
      RECT 1.000000 44.430000 40.020000 45.040000 ;
      RECT 0.000000 44.190000 40.020000 44.430000 ;
      RECT 1.000000 43.720000 40.020000 44.190000 ;
      RECT 1.000000 43.210000 2.530000 43.720000 ;
      RECT 0.000000 42.970000 2.530000 43.210000 ;
      RECT 37.490000 42.640000 40.020000 43.720000 ;
      RECT 8.560000 42.640000 35.690000 43.720000 ;
      RECT 4.330000 42.640000 6.760000 43.720000 ;
      RECT 1.000000 42.640000 2.530000 42.970000 ;
      RECT 1.000000 42.360000 40.020000 42.640000 ;
      RECT 1.000000 41.990000 39.020000 42.360000 ;
      RECT 0.000000 41.380000 39.020000 41.990000 ;
      RECT 0.000000 41.140000 40.020000 41.380000 ;
      RECT 1.000000 41.000000 40.020000 41.140000 ;
      RECT 39.290000 39.920000 40.020000 41.000000 ;
      RECT 6.560000 39.920000 37.490000 41.000000 ;
      RECT 2.530000 39.920000 4.595000 41.000000 ;
      RECT 0.000000 39.920000 0.730000 40.160000 ;
      RECT 1.000000 38.940000 40.020000 39.920000 ;
      RECT 0.000000 38.700000 40.020000 38.940000 ;
      RECT 0.000000 38.280000 39.020000 38.700000 ;
      RECT 0.000000 38.090000 2.530000 38.280000 ;
      RECT 37.490000 37.720000 39.020000 38.280000 ;
      RECT 37.490000 37.200000 40.020000 37.720000 ;
      RECT 8.560000 37.200000 35.690000 38.280000 ;
      RECT 4.330000 37.200000 6.760000 38.280000 ;
      RECT 1.000000 37.200000 2.530000 38.090000 ;
      RECT 1.000000 37.110000 40.020000 37.200000 ;
      RECT 0.000000 36.870000 40.020000 37.110000 ;
      RECT 1.000000 35.890000 40.020000 36.870000 ;
      RECT 0.000000 35.560000 40.020000 35.890000 ;
      RECT 39.290000 35.040000 40.020000 35.560000 ;
      RECT 0.000000 35.040000 0.730000 35.560000 ;
      RECT 6.560000 34.480000 37.490000 35.560000 ;
      RECT 2.530000 34.480000 4.595000 35.560000 ;
      RECT 1.000000 34.060000 39.020000 34.480000 ;
      RECT 0.000000 33.820000 40.020000 34.060000 ;
      RECT 1.000000 32.840000 40.020000 33.820000 ;
      RECT 0.000000 31.990000 2.530000 32.840000 ;
      RECT 37.490000 31.760000 40.020000 32.840000 ;
      RECT 8.560000 31.760000 35.690000 32.840000 ;
      RECT 4.330000 31.760000 6.760000 32.840000 ;
      RECT 1.000000 31.760000 2.530000 31.990000 ;
      RECT 1.000000 31.380000 40.020000 31.760000 ;
      RECT 1.000000 31.010000 39.020000 31.380000 ;
      RECT 0.000000 30.770000 39.020000 31.010000 ;
      RECT 1.000000 30.400000 39.020000 30.770000 ;
      RECT 1.000000 30.120000 40.020000 30.400000 ;
      RECT 0.000000 29.550000 0.730000 29.790000 ;
      RECT 39.290000 29.040000 40.020000 30.120000 ;
      RECT 6.560000 29.040000 37.490000 30.120000 ;
      RECT 2.530000 29.040000 4.595000 30.120000 ;
      RECT 1.000000 28.570000 40.020000 29.040000 ;
      RECT 0.000000 27.720000 40.020000 28.570000 ;
      RECT 1.000000 27.400000 39.020000 27.720000 ;
      RECT 37.490000 26.740000 39.020000 27.400000 ;
      RECT 1.000000 26.740000 2.530000 27.400000 ;
      RECT 0.000000 26.500000 2.530000 26.740000 ;
      RECT 37.490000 26.320000 40.020000 26.740000 ;
      RECT 8.560000 26.320000 35.690000 27.400000 ;
      RECT 4.330000 26.320000 6.760000 27.400000 ;
      RECT 1.000000 26.320000 2.530000 26.500000 ;
      RECT 1.000000 25.520000 40.020000 26.320000 ;
      RECT 0.000000 24.680000 40.020000 25.520000 ;
      RECT 0.000000 24.670000 0.730000 24.680000 ;
      RECT 39.290000 24.060000 40.020000 24.680000 ;
      RECT 6.560000 23.600000 37.490000 24.680000 ;
      RECT 2.530000 23.600000 4.595000 24.680000 ;
      RECT 0.000000 23.600000 0.730000 23.690000 ;
      RECT 0.000000 23.450000 39.020000 23.600000 ;
      RECT 1.000000 23.080000 39.020000 23.450000 ;
      RECT 1.000000 22.470000 40.020000 23.080000 ;
      RECT 0.000000 21.960000 40.020000 22.470000 ;
      RECT 0.000000 21.620000 2.530000 21.960000 ;
      RECT 37.490000 20.880000 40.020000 21.960000 ;
      RECT 8.560000 20.880000 35.690000 21.960000 ;
      RECT 4.330000 20.880000 6.760000 21.960000 ;
      RECT 1.000000 20.880000 2.530000 21.620000 ;
      RECT 1.000000 20.640000 40.020000 20.880000 ;
      RECT 0.000000 20.400000 40.020000 20.640000 ;
      RECT 1.000000 19.420000 39.020000 20.400000 ;
      RECT 0.000000 19.240000 40.020000 19.420000 ;
      RECT 0.000000 18.570000 0.730000 19.240000 ;
      RECT 39.290000 18.160000 40.020000 19.240000 ;
      RECT 6.560000 18.160000 37.490000 19.240000 ;
      RECT 2.530000 18.160000 4.595000 19.240000 ;
      RECT 1.000000 17.590000 40.020000 18.160000 ;
      RECT 0.000000 17.350000 40.020000 17.590000 ;
      RECT 1.000000 16.740000 40.020000 17.350000 ;
      RECT 1.000000 16.520000 39.020000 16.740000 ;
      RECT 1.000000 16.370000 2.530000 16.520000 ;
      RECT 0.000000 16.130000 2.530000 16.370000 ;
      RECT 37.490000 15.760000 39.020000 16.520000 ;
      RECT 37.490000 15.440000 40.020000 15.760000 ;
      RECT 8.560000 15.440000 35.690000 16.520000 ;
      RECT 4.330000 15.440000 6.760000 16.520000 ;
      RECT 1.000000 15.440000 2.530000 16.130000 ;
      RECT 1.000000 15.150000 40.020000 15.440000 ;
      RECT 0.000000 14.300000 40.020000 15.150000 ;
      RECT 1.000000 13.800000 40.020000 14.300000 ;
      RECT 39.290000 13.080000 40.020000 13.800000 ;
      RECT 0.000000 13.080000 0.730000 13.320000 ;
      RECT 6.560000 12.720000 37.490000 13.800000 ;
      RECT 2.530000 12.720000 4.595000 13.800000 ;
      RECT 1.000000 12.100000 39.020000 12.720000 ;
      RECT 0.000000 11.250000 40.020000 12.100000 ;
      RECT 1.000000 11.080000 40.020000 11.250000 ;
      RECT 1.000000 10.270000 2.530000 11.080000 ;
      RECT 0.000000 10.030000 2.530000 10.270000 ;
      RECT 37.490000 10.000000 40.020000 11.080000 ;
      RECT 8.560000 10.000000 35.690000 11.080000 ;
      RECT 4.330000 10.000000 6.760000 11.080000 ;
      RECT 1.000000 10.000000 2.530000 10.030000 ;
      RECT 1.000000 9.420000 40.020000 10.000000 ;
      RECT 1.000000 9.050000 39.020000 9.420000 ;
      RECT 0.000000 8.440000 39.020000 9.050000 ;
      RECT 0.000000 8.360000 40.020000 8.440000 ;
      RECT 0.000000 8.200000 0.730000 8.360000 ;
      RECT 39.290000 7.280000 40.020000 8.360000 ;
      RECT 6.560000 7.280000 37.490000 8.360000 ;
      RECT 2.530000 7.280000 4.595000 8.360000 ;
      RECT 1.000000 7.220000 40.020000 7.280000 ;
      RECT 0.000000 6.980000 40.020000 7.220000 ;
      RECT 1.000000 6.000000 40.020000 6.980000 ;
      RECT 0.000000 5.760000 40.020000 6.000000 ;
      RECT 1.000000 5.640000 39.020000 5.760000 ;
      RECT 37.490000 4.780000 39.020000 5.640000 ;
      RECT 1.000000 4.780000 2.530000 5.640000 ;
      RECT 37.490000 4.560000 40.020000 4.780000 ;
      RECT 8.560000 4.560000 35.690000 5.640000 ;
      RECT 4.330000 4.560000 6.760000 5.640000 ;
      RECT 0.000000 4.560000 2.530000 4.780000 ;
      RECT 0.000000 4.350000 40.020000 4.560000 ;
      RECT 0.000000 0.000000 40.020000 0.750000 ;
    LAYER met4 ;
      RECT 4.330000 198.320000 35.690000 200.260000 ;
      RECT 6.560000 196.520000 35.690000 198.320000 ;
      RECT 4.330000 193.320000 4.760000 198.320000 ;
      RECT 4.330000 192.240000 4.595000 193.320000 ;
      RECT 4.330000 187.880000 4.760000 192.240000 ;
      RECT 4.330000 186.800000 4.595000 187.880000 ;
      RECT 4.330000 182.440000 4.760000 186.800000 ;
      RECT 4.330000 181.360000 4.595000 182.440000 ;
      RECT 4.330000 177.000000 4.760000 181.360000 ;
      RECT 4.330000 175.920000 4.595000 177.000000 ;
      RECT 4.330000 171.560000 4.760000 175.920000 ;
      RECT 4.330000 170.480000 4.595000 171.560000 ;
      RECT 4.330000 166.120000 4.760000 170.480000 ;
      RECT 4.330000 165.040000 4.595000 166.120000 ;
      RECT 4.330000 160.680000 4.760000 165.040000 ;
      RECT 4.330000 159.600000 4.595000 160.680000 ;
      RECT 4.330000 155.240000 4.760000 159.600000 ;
      RECT 4.330000 154.160000 4.595000 155.240000 ;
      RECT 4.330000 149.800000 4.760000 154.160000 ;
      RECT 4.330000 148.720000 4.595000 149.800000 ;
      RECT 4.330000 144.360000 4.760000 148.720000 ;
      RECT 4.330000 143.280000 4.595000 144.360000 ;
      RECT 4.330000 138.920000 4.760000 143.280000 ;
      RECT 4.330000 137.840000 4.595000 138.920000 ;
      RECT 4.330000 133.480000 4.760000 137.840000 ;
      RECT 4.330000 132.400000 4.595000 133.480000 ;
      RECT 4.330000 128.040000 4.760000 132.400000 ;
      RECT 4.330000 126.960000 4.595000 128.040000 ;
      RECT 4.330000 122.600000 4.760000 126.960000 ;
      RECT 4.330000 121.520000 4.595000 122.600000 ;
      RECT 4.330000 117.160000 4.760000 121.520000 ;
      RECT 4.330000 116.080000 4.595000 117.160000 ;
      RECT 4.330000 111.720000 4.760000 116.080000 ;
      RECT 4.330000 110.640000 4.595000 111.720000 ;
      RECT 4.330000 106.280000 4.760000 110.640000 ;
      RECT 4.330000 105.200000 4.595000 106.280000 ;
      RECT 4.330000 100.840000 4.760000 105.200000 ;
      RECT 4.330000 99.760000 4.595000 100.840000 ;
      RECT 4.330000 95.400000 4.760000 99.760000 ;
      RECT 4.330000 94.320000 4.595000 95.400000 ;
      RECT 4.330000 89.960000 4.760000 94.320000 ;
      RECT 4.330000 88.880000 4.595000 89.960000 ;
      RECT 4.330000 84.520000 4.760000 88.880000 ;
      RECT 4.330000 83.440000 4.595000 84.520000 ;
      RECT 4.330000 79.080000 4.760000 83.440000 ;
      RECT 4.330000 78.000000 4.595000 79.080000 ;
      RECT 4.330000 73.640000 4.760000 78.000000 ;
      RECT 4.330000 72.560000 4.595000 73.640000 ;
      RECT 4.330000 68.200000 4.760000 72.560000 ;
      RECT 4.330000 67.120000 4.595000 68.200000 ;
      RECT 4.330000 62.760000 4.760000 67.120000 ;
      RECT 4.330000 61.680000 4.595000 62.760000 ;
      RECT 4.330000 57.320000 4.760000 61.680000 ;
      RECT 4.330000 56.240000 4.595000 57.320000 ;
      RECT 4.330000 51.880000 4.760000 56.240000 ;
      RECT 4.330000 50.800000 4.595000 51.880000 ;
      RECT 4.330000 46.440000 4.760000 50.800000 ;
      RECT 4.330000 45.360000 4.595000 46.440000 ;
      RECT 4.330000 41.000000 4.760000 45.360000 ;
      RECT 4.330000 39.920000 4.595000 41.000000 ;
      RECT 4.330000 35.560000 4.760000 39.920000 ;
      RECT 4.330000 34.480000 4.595000 35.560000 ;
      RECT 4.330000 30.120000 4.760000 34.480000 ;
      RECT 4.330000 29.040000 4.595000 30.120000 ;
      RECT 4.330000 24.680000 4.760000 29.040000 ;
      RECT 4.330000 23.600000 4.595000 24.680000 ;
      RECT 4.330000 19.240000 4.760000 23.600000 ;
      RECT 4.330000 18.160000 4.595000 19.240000 ;
      RECT 4.330000 13.800000 4.760000 18.160000 ;
      RECT 4.330000 12.720000 4.595000 13.800000 ;
      RECT 4.330000 8.360000 4.760000 12.720000 ;
      RECT 4.330000 7.280000 4.595000 8.360000 ;
      RECT 8.560000 2.550000 35.690000 196.520000 ;
      RECT 6.560000 2.550000 6.760000 196.520000 ;
      RECT 6.560000 0.750000 35.690000 2.550000 ;
      RECT 4.330000 0.750000 4.760000 7.280000 ;
      RECT 39.290000 0.000000 40.020000 200.260000 ;
      RECT 4.330000 0.000000 35.690000 0.750000 ;
      RECT 0.000000 0.000000 0.730000 200.260000 ;
  END
END E_CPU_IO

END LIBRARY
