##
## LEF for PtnCells ;
## created by Innovus v19.11-s128_1 on Wed Dec  8 10:37:29 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO BlockRAM_1KB
  CLASS BLOCK ;
  SIZE 529.920000 BY 420.240000 ;
  FOREIGN BlockRAM_1KB 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5773 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.0457 LAYER met3  ;
    ANTENNAMAXAREACAR 23.1899 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 107.705 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.488562 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 63.7624 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 341.304 LAYER met4  ;
    ANTENNAGATEAREA 5.8407 LAYER met4  ;
    ANTENNAMAXAREACAR 91.7241 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 459.439 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.524528 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 200.280000 0.720000 200.660000 ;
    END
  END clk
  PIN rd_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.6467 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 110.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 53.7361 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 267.297 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6602 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.672 LAYER met4  ;
    ANTENNAGATEAREA 0.4347 LAYER met4  ;
    ANTENNAMAXAREACAR 55.2549 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 275.744 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 85.600000 0.720000 85.980000 ;
    END
  END rd_addr[7]
  PIN rd_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.3135 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 93.896 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met4  ;
    ANTENNAMAXAREACAR 46.7582 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 233.6 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 88.650000 0.720000 89.030000 ;
    END
  END rd_addr[6]
  PIN rd_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.7324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.368 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 71.8979 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 349.013 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.8562 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.384 LAYER met4  ;
    ANTENNAGATEAREA 0.4347 LAYER met4  ;
    ANTENNAMAXAREACAR 78.4684 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 384.403 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 92.310000 0.720000 92.690000 ;
    END
  END rd_addr[5]
  PIN rd_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.1324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.168 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 84.608 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 407.167 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.5562 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.784 LAYER met4  ;
    ANTENNAGATEAREA 0.4347 LAYER met4  ;
    ANTENNAMAXAREACAR 90.4884 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 438.876 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 95.360000 0.720000 95.740000 ;
    END
  END rd_addr[4]
  PIN rd_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.4464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.664 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 22.6655 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 98.1493 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 72.180000 0.720000 72.560000 ;
    END
  END rd_addr[3]
  PIN rd_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 75.3944 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 402.72 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 202.329 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1052.06 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 75.230000 0.720000 75.610000 ;
    END
  END rd_addr[2]
  PIN rd_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.2994 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.392 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.4444 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 206.448 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met4  ;
    ANTENNAMAXAREACAR 100.607 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 520.097 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 78.890000 0.720000 79.270000 ;
    END
  END rd_addr[1]
  PIN rd_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.1434 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.56 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 202.387 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 991.613 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.512537 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.8782 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.168 LAYER met4  ;
    ANTENNAGATEAREA 0.4347 LAYER met4  ;
    ANTENNAMAXAREACAR 206.708 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1015 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.512537 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 81.940000 0.720000 82.320000 ;
    END
  END rd_addr[0]
  PIN rd_data[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.7592 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.848 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 261.890000 0.720000 262.270000 ;
    END
  END rd_data[31]
  PIN rd_data[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6594 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.2788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 204.624 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 266.770000 0.720000 267.150000 ;
    END
  END rd_data[30]
  PIN rd_data[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.472 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 271.040000 0.720000 271.420000 ;
    END
  END rd_data[29]
  PIN rd_data[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.4258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.408 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 275.920000 0.720000 276.300000 ;
    END
  END rd_data[28]
  PIN rd_data[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7294 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 61.9464 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 331.792 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 242.980000 0.720000 243.360000 ;
    END
  END rd_data[27]
  PIN rd_data[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.2272 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 247.860000 0.720000 248.240000 ;
    END
  END rd_data[26]
  PIN rd_data[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.4144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 252.130000 0.720000 252.510000 ;
    END
  END rd_data[25]
  PIN rd_data[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.992 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 257.010000 0.720000 257.390000 ;
    END
  END rd_data[24]
  PIN rd_data[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.736 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 224.070000 0.720000 224.450000 ;
    END
  END rd_data[23]
  PIN rd_data[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.4258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.408 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 228.340000 0.720000 228.720000 ;
    END
  END rd_data[22]
  PIN rd_data[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.472 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 233.220000 0.720000 233.600000 ;
    END
  END rd_data[21]
  PIN rd_data[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.208 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 238.100000 0.720000 238.480000 ;
    END
  END rd_data[20]
  PIN rd_data[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5544 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.2428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.432 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 205.160000 0.720000 205.540000 ;
    END
  END rd_data[19]
  PIN rd_data[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5414 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.216 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 209.430000 0.720000 209.810000 ;
    END
  END rd_data[18]
  PIN rd_data[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5754 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.064 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 214.310000 0.720000 214.690000 ;
    END
  END rd_data[17]
  PIN rd_data[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4546 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.3568 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 253.04 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 219.190000 0.720000 219.570000 ;
    END
  END rd_data[16]
  PIN rd_data[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.5008 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.808 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 45.340000 0.720000 45.720000 ;
    END
  END rd_data[15]
  PIN rd_data[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.9814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.896 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 48.390000 0.720000 48.770000 ;
    END
  END rd_data[14]
  PIN rd_data[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.1904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 52.050000 0.720000 52.430000 ;
    END
  END rd_data[13]
  PIN rd_data[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.1224 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.648 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 55.100000 0.720000 55.480000 ;
    END
  END rd_data[12]
  PIN rd_data[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5216 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.8688 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 245.104 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 31.920000 0.720000 32.300000 ;
    END
  END rd_data[11]
  PIN rd_data[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9036 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 80.1378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 427.872 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 34.970000 0.720000 35.350000 ;
    END
  END rd_data[10]
  PIN rd_data[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.6808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.768 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 38.630000 0.720000 39.010000 ;
    END
  END rd_data[9]
  PIN rd_data[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.472 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 41.680000 0.720000 42.060000 ;
    END
  END rd_data[8]
  PIN rd_data[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4436 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.024 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.1578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.312 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 18.500000 0.720000 18.880000 ;
    END
  END rd_data[7]
  PIN rd_data[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6186 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 64.2966 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 343.856 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 21.550000 0.720000 21.930000 ;
    END
  END rd_data[6]
  PIN rd_data[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.208 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 25.210000 0.720000 25.590000 ;
    END
  END rd_data[5]
  PIN rd_data[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8956 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.2496 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 162.272 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 28.260000 0.720000 28.640000 ;
    END
  END rd_data[4]
  PIN rd_data[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.472 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 5.080000 0.720000 5.460000 ;
    END
  END rd_data[3]
  PIN rd_data[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8686 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 98.5098 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 525.856 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 8.130000 0.720000 8.510000 ;
    END
  END rd_data[2]
  PIN rd_data[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4706 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 110.111 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 587.728 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 11.790000 0.720000 12.170000 ;
    END
  END rd_data[1]
  PIN rd_data[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 14.840000 0.720000 15.220000 ;
    END
  END rd_data[0]
  PIN wr_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.7256 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 68.2763 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 330.385 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 309.470000 0.720000 309.850000 ;
    END
  END wr_addr[7]
  PIN wr_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.2056 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 68.3009 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 328.622 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 313.740000 0.720000 314.120000 ;
    END
  END wr_addr[6]
  PIN wr_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.7068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 36.24 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met4  ;
    ANTENNAMAXAREACAR 81.7088 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 403.343 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 318.620000 0.720000 319.000000 ;
    END
  END wr_addr[5]
  PIN wr_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.7216 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.328 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 83.1822 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 405.407 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 323.500000 0.720000 323.880000 ;
    END
  END wr_addr[4]
  PIN wr_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.6496 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 78.7062 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 383.389 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 290.560000 0.720000 290.940000 ;
    END
  END wr_addr[3]
  PIN wr_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.4466 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.528 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 73.6959 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 357.325 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 294.830000 0.720000 295.210000 ;
    END
  END wr_addr[2]
  PIN wr_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.8526 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.872 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.2076 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 258.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met4  ;
    ANTENNAMAXAREACAR 127.177 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 658.045 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 299.710000 0.720000 300.090000 ;
    END
  END wr_addr[1]
  PIN wr_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6326 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 88.616 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 473.24 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met4  ;
    ANTENNAMAXAREACAR 225.896 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1185.46 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.486312 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 304.590000 0.720000 304.970000 ;
    END
  END wr_addr[0]
  PIN wr_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.6182 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.096 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met3  ;
    ANTENNAMAXAREACAR 38.9834 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 182.116 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.479276 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 385.110000 0.720000 385.490000 ;
    END
  END wr_data[31]
  PIN wr_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5756 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 121.69 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 649.952 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 358.118 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1849.15 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.550615 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 389.990000 0.720000 390.370000 ;
    END
  END wr_data[30]
  PIN wr_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9896 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 77.1858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 412.128 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 194.962 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1005.38 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.729187 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 394.870000 0.720000 395.250000 ;
    END
  END wr_data[29]
  PIN wr_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 117.016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 625.024 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 289.847 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1522 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.729187 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 399.140000 0.720000 399.520000 ;
    END
  END wr_data[28]
  PIN wr_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met3  ;
    ANTENNAMAXAREACAR 116.72 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 564.903 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.479276 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 366.200000 0.720000 366.580000 ;
    END
  END wr_data[27]
  PIN wr_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.8204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.704 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met3  ;
    ANTENNAMAXAREACAR 117.86 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 575.453 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.479276 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 371.080000 0.720000 371.460000 ;
    END
  END wr_data[26]
  PIN wr_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1616 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 303.664 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met4  ;
    ANTENNAMAXAREACAR 117.465 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 606.867 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.703007 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 375.960000 0.720000 376.340000 ;
    END
  END wr_data[25]
  PIN wr_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8716 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 61.1298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 326.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met4  ;
    ANTENNAMAXAREACAR 129.839 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 662.138 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.524436 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 380.230000 0.720000 380.610000 ;
    END
  END wr_data[24]
  PIN wr_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4116 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.6578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 217.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 123.373 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 626.609 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.412172 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 347.290000 0.720000 347.670000 ;
    END
  END wr_data[23]
  PIN wr_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 91.6428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 489.232 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 185.892 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 970.282 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.550615 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 352.170000 0.720000 352.550000 ;
    END
  END wr_data[22]
  PIN wr_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.8726 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 506.928 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 179.558 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 938.323 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.550615 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 356.440000 0.720000 356.820000 ;
    END
  END wr_data[21]
  PIN wr_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.0326 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 92.9958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 496.448 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0557 LAYER met4  ;
    ANTENNAMAXAREACAR 101.361 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 520.694 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.483716 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 361.320000 0.720000 361.700000 ;
    END
  END wr_data[20]
  PIN wr_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.3042 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.088 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met3  ;
    ANTENNAMAXAREACAR 23.562 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 104.113 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.479276 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 328.380000 0.720000 328.760000 ;
    END
  END wr_data[19]
  PIN wr_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.9286 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 83.0418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 443.36 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 180.369 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 937.47 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.550615 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 333.260000 0.720000 333.640000 ;
    END
  END wr_data[18]
  PIN wr_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6426 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.8558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 250.368 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1717 LAYER met4  ;
    ANTENNAMAXAREACAR 37.2516 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 176.274 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.444774 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 337.530000 0.720000 337.910000 ;
    END
  END wr_data[17]
  PIN wr_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2856 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 71.4888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 381.744 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9287 LAYER met4  ;
    ANTENNAMAXAREACAR 46.6687 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 229.621 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.449415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 342.410000 0.720000 342.790000 ;
    END
  END wr_data[16]
  PIN wr_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.0184 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.76 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 38.9975 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 178.189 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.874123 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 139.280000 0.720000 139.660000 ;
    END
  END wr_data[15]
  PIN wr_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.9344 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 32.617 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 145.819 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.466186 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 142.330000 0.720000 142.710000 ;
    END
  END wr_data[14]
  PIN wr_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8256 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.4766 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 104.816 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met4  ;
    ANTENNAMAXAREACAR 46.3846 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 225.571 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.524436 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 145.990000 0.720000 146.370000 ;
    END
  END wr_data[13]
  PIN wr_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.9914 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.616 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 37.2024 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 170.072 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.466186 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 149.040000 0.720000 149.420000 ;
    END
  END wr_data[12]
  PIN wr_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.0164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 44.7634 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 73.1134 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.466186 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 125.860000 0.720000 126.240000 ;
    END
  END wr_data[11]
  PIN wr_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1544 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.152 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 32.2155 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 143.111 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.644758 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 128.910000 0.720000 129.290000 ;
    END
  END wr_data[10]
  PIN wr_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.5074 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.368 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 21.6586 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 91.1618 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.466186 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 132.570000 0.720000 132.950000 ;
    END
  END wr_data[9]
  PIN wr_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.736 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 18.7437 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 75.0564 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.644758 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 135.620000 0.720000 136.000000 ;
    END
  END wr_data[8]
  PIN wr_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.2124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.928 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 42.4091 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 203.67 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.761257 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.4028 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 83.24 LAYER met4  ;
    ANTENNAGATEAREA 0.6867 LAYER met4  ;
    ANTENNAMAXAREACAR 64.8393 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 324.888 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.761257 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 112.440000 0.720000 112.820000 ;
    END
  END wr_data[7]
  PIN wr_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 49.7614 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 265.856 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 107.699 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 551.153 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.761257 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.1812 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.784 LAYER met4  ;
    ANTENNAGATEAREA 0.6867 LAYER met4  ;
    ANTENNAMAXAREACAR 110.876 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 568.314 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.761257 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 115.490000 0.720000 115.870000 ;
    END
  END wr_data[6]
  PIN wr_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.0608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 129.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met4  ;
    ANTENNAMAXAREACAR 110.953 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 577.983 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.640935 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 119.150000 0.720000 119.530000 ;
    END
  END wr_data[5]
  PIN wr_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.7944 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.032 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 48.837 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 231.833 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.582685 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.834 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 111.736 LAYER met4  ;
    ANTENNAGATEAREA 0.6867 LAYER met4  ;
    ANTENNAMAXAREACAR 79.1763 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 394.547 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.582685 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 122.200000 0.720000 122.580000 ;
    END
  END wr_data[4]
  PIN wr_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.3512 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.472 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 31.5521 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 142.865 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.582685 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5212 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.264 LAYER met4  ;
    ANTENNAGATEAREA 0.6867 LAYER met4  ;
    ANTENNAMAXAREACAR 33.7674 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 154.899 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.582685 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 99.020000 0.720000 99.400000 ;
    END
  END wr_data[3]
  PIN wr_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2636 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.188 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 97.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met4  ;
    ANTENNAMAXAREACAR 51.7395 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 257.774 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.640935 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 102.070000 0.720000 102.450000 ;
    END
  END wr_data[2]
  PIN wr_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.304 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met3  ;
    ANTENNAMAXAREACAR 39.5339 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 188.003 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.582685 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5752 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.552 LAYER met4  ;
    ANTENNAGATEAREA 0.6867 LAYER met4  ;
    ANTENNAMAXAREACAR 41.8278 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 200.457 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.582685 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 105.730000 0.720000 106.110000 ;
    END
  END wr_data[1]
  PIN wr_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.8578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 123 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6867 LAYER met4  ;
    ANTENNAMAXAREACAR 43.7865 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 218.846 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.640935 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 108.780000 0.720000 109.160000 ;
    END
  END wr_data[0]
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.0864 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.456 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0457 LAYER met3  ;
    ANTENNAMAXAREACAR 8.73208 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 35.5795 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.28515 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 68.520000 0.720000 68.900000 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.0864 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.456 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6767 LAYER met3  ;
    ANTENNAMAXAREACAR 11.9922 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 49.7212 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.431793 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 65.470000 0.720000 65.850000 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6156 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.0858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.928 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.4247 LAYER met4  ;
    ANTENNAMAXAREACAR 22.2522 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 99.1785 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.130329 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 61.810000 0.720000 62.190000 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1796 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.9296 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 139.232 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1817 LAYER met4  ;
    ANTENNAMAXAREACAR 29.5126 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 147.298 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.654207 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 58.760000 0.720000 59.140000 ;
    END
  END C3
  PIN C4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6266 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 62.5938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 334.304 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9297 LAYER met4  ;
    ANTENNAMAXAREACAR 75.6987 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 383.989 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.204292 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 285.680000 0.720000 286.060000 ;
    END
  END C4
  PIN C5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.344 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 8.4987 LAYER met3  ;
    ANTENNAMAXAREACAR 15.5497 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 64.7059 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.308054 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 280.800000 0.720000 281.180000 ;
    END
  END C5
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 529.120000 415.570000 529.920000 416.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 529.120000 2.850000 529.920000 3.650000 ;
    END
    PORT
      LAYER met4 ;
        RECT 526.290000 419.440000 527.090000 420.240000 ;
    END
    PORT
      LAYER met4 ;
        RECT 526.290000 0.000000 527.090000 0.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 419.440000 3.630000 420.240000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 0.000000 3.630000 0.800000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 2.830000 2.850000 529.920000 3.650000 ;
        RECT 2.830000 415.570000 529.920000 416.370000 ;
        RECT 2.830000 10.300000 3.630000 10.780000 ;
        RECT 2.830000 4.860000 3.630000 5.340000 ;
        RECT 2.830000 15.740000 3.630000 16.220000 ;
        RECT 2.830000 21.180000 3.630000 21.660000 ;
        RECT 2.830000 26.620000 3.630000 27.100000 ;
        RECT 2.830000 32.060000 3.630000 32.540000 ;
        RECT 2.830000 37.500000 3.630000 37.980000 ;
        RECT 2.830000 42.940000 3.630000 43.420000 ;
        RECT 2.830000 48.380000 3.630000 48.860000 ;
        RECT 2.830000 53.820000 3.630000 54.300000 ;
        RECT 2.830000 59.260000 3.630000 59.740000 ;
        RECT 2.830000 64.700000 3.630000 65.180000 ;
        RECT 2.830000 70.140000 3.630000 70.620000 ;
        RECT 2.830000 75.580000 3.630000 76.060000 ;
        RECT 2.830000 81.020000 3.630000 81.500000 ;
        RECT 2.830000 86.460000 3.630000 86.940000 ;
        RECT 2.830000 91.900000 3.630000 92.380000 ;
        RECT 2.830000 97.340000 3.630000 97.820000 ;
        RECT 2.830000 102.780000 3.630000 103.260000 ;
        RECT 2.830000 108.220000 3.630000 108.700000 ;
        RECT 2.830000 113.660000 3.630000 114.140000 ;
        RECT 2.830000 119.100000 3.630000 119.580000 ;
        RECT 2.830000 124.540000 3.630000 125.020000 ;
        RECT 2.830000 140.860000 3.630000 141.340000 ;
        RECT 2.830000 135.420000 3.630000 135.900000 ;
        RECT 2.830000 129.980000 3.630000 130.460000 ;
        RECT 2.830000 146.300000 3.630000 146.780000 ;
        RECT 2.830000 151.740000 3.630000 152.220000 ;
        RECT 2.830000 157.180000 3.630000 157.660000 ;
        RECT 2.830000 162.620000 3.630000 163.100000 ;
        RECT 2.830000 168.060000 3.630000 168.540000 ;
        RECT 2.830000 173.500000 3.630000 173.980000 ;
        RECT 2.830000 178.940000 3.630000 179.420000 ;
        RECT 2.830000 184.380000 3.630000 184.860000 ;
        RECT 2.830000 189.820000 3.630000 190.300000 ;
        RECT 2.830000 195.260000 3.630000 195.740000 ;
        RECT 2.830000 200.700000 3.630000 201.180000 ;
        RECT 2.830000 206.140000 3.630000 206.620000 ;
        RECT 526.290000 10.300000 527.090000 10.780000 ;
        RECT 526.290000 4.860000 527.090000 5.340000 ;
        RECT 526.290000 15.740000 527.090000 16.220000 ;
        RECT 526.290000 21.180000 527.090000 21.660000 ;
        RECT 526.290000 26.620000 527.090000 27.100000 ;
        RECT 526.290000 32.060000 527.090000 32.540000 ;
        RECT 526.290000 37.500000 527.090000 37.980000 ;
        RECT 526.290000 42.940000 527.090000 43.420000 ;
        RECT 526.290000 48.380000 527.090000 48.860000 ;
        RECT 526.290000 53.820000 527.090000 54.300000 ;
        RECT 526.290000 59.260000 527.090000 59.740000 ;
        RECT 526.290000 64.700000 527.090000 65.180000 ;
        RECT 526.290000 70.140000 527.090000 70.620000 ;
        RECT 526.290000 75.580000 527.090000 76.060000 ;
        RECT 526.290000 81.020000 527.090000 81.500000 ;
        RECT 526.290000 86.460000 527.090000 86.940000 ;
        RECT 526.290000 91.900000 527.090000 92.380000 ;
        RECT 526.290000 97.340000 527.090000 97.820000 ;
        RECT 526.290000 102.780000 527.090000 103.260000 ;
        RECT 526.290000 108.220000 527.090000 108.700000 ;
        RECT 526.290000 113.660000 527.090000 114.140000 ;
        RECT 526.290000 119.100000 527.090000 119.580000 ;
        RECT 526.290000 124.540000 527.090000 125.020000 ;
        RECT 526.290000 140.860000 527.090000 141.340000 ;
        RECT 526.290000 135.420000 527.090000 135.900000 ;
        RECT 526.290000 129.980000 527.090000 130.460000 ;
        RECT 526.290000 146.300000 527.090000 146.780000 ;
        RECT 526.290000 151.740000 527.090000 152.220000 ;
        RECT 526.290000 157.180000 527.090000 157.660000 ;
        RECT 526.290000 162.620000 527.090000 163.100000 ;
        RECT 526.290000 168.060000 527.090000 168.540000 ;
        RECT 526.290000 173.500000 527.090000 173.980000 ;
        RECT 526.290000 178.940000 527.090000 179.420000 ;
        RECT 526.290000 184.380000 527.090000 184.860000 ;
        RECT 526.290000 189.820000 527.090000 190.300000 ;
        RECT 526.290000 195.260000 527.090000 195.740000 ;
        RECT 526.290000 200.700000 527.090000 201.180000 ;
        RECT 526.290000 206.140000 527.090000 206.620000 ;
        RECT 2.830000 342.140000 3.630000 342.620000 ;
        RECT 2.830000 211.580000 3.630000 212.060000 ;
        RECT 2.830000 217.020000 3.630000 217.500000 ;
        RECT 2.830000 222.460000 3.630000 222.940000 ;
        RECT 2.830000 227.900000 3.630000 228.380000 ;
        RECT 2.830000 233.340000 3.630000 233.820000 ;
        RECT 2.830000 238.780000 3.630000 239.260000 ;
        RECT 2.830000 244.220000 3.630000 244.700000 ;
        RECT 2.830000 249.660000 3.630000 250.140000 ;
        RECT 2.830000 255.100000 3.630000 255.580000 ;
        RECT 2.830000 260.540000 3.630000 261.020000 ;
        RECT 2.830000 265.980000 3.630000 266.460000 ;
        RECT 2.830000 271.420000 3.630000 271.900000 ;
        RECT 2.830000 276.860000 3.630000 277.340000 ;
        RECT 2.830000 282.300000 3.630000 282.780000 ;
        RECT 2.830000 287.740000 3.630000 288.220000 ;
        RECT 2.830000 293.180000 3.630000 293.660000 ;
        RECT 2.830000 298.620000 3.630000 299.100000 ;
        RECT 2.830000 304.060000 3.630000 304.540000 ;
        RECT 2.830000 325.820000 3.630000 326.300000 ;
        RECT 2.830000 309.500000 3.630000 309.980000 ;
        RECT 2.830000 314.940000 3.630000 315.420000 ;
        RECT 2.830000 320.380000 3.630000 320.860000 ;
        RECT 2.830000 336.700000 3.630000 337.180000 ;
        RECT 2.830000 331.260000 3.630000 331.740000 ;
        RECT 2.830000 347.580000 3.630000 348.060000 ;
        RECT 2.830000 353.020000 3.630000 353.500000 ;
        RECT 2.830000 358.460000 3.630000 358.940000 ;
        RECT 2.830000 363.900000 3.630000 364.380000 ;
        RECT 2.830000 369.340000 3.630000 369.820000 ;
        RECT 2.830000 374.780000 3.630000 375.260000 ;
        RECT 2.830000 380.220000 3.630000 380.700000 ;
        RECT 2.830000 385.660000 3.630000 386.140000 ;
        RECT 2.830000 391.100000 3.630000 391.580000 ;
        RECT 2.830000 396.540000 3.630000 397.020000 ;
        RECT 2.830000 401.980000 3.630000 402.460000 ;
        RECT 2.830000 407.420000 3.630000 407.900000 ;
        RECT 2.830000 412.860000 3.630000 413.340000 ;
        RECT 526.290000 342.140000 527.090000 342.620000 ;
        RECT 526.290000 211.580000 527.090000 212.060000 ;
        RECT 526.290000 217.020000 527.090000 217.500000 ;
        RECT 526.290000 222.460000 527.090000 222.940000 ;
        RECT 526.290000 227.900000 527.090000 228.380000 ;
        RECT 526.290000 233.340000 527.090000 233.820000 ;
        RECT 526.290000 238.780000 527.090000 239.260000 ;
        RECT 526.290000 244.220000 527.090000 244.700000 ;
        RECT 526.290000 249.660000 527.090000 250.140000 ;
        RECT 526.290000 255.100000 527.090000 255.580000 ;
        RECT 526.290000 260.540000 527.090000 261.020000 ;
        RECT 526.290000 265.980000 527.090000 266.460000 ;
        RECT 526.290000 271.420000 527.090000 271.900000 ;
        RECT 526.290000 276.860000 527.090000 277.340000 ;
        RECT 526.290000 282.300000 527.090000 282.780000 ;
        RECT 526.290000 287.740000 527.090000 288.220000 ;
        RECT 526.290000 293.180000 527.090000 293.660000 ;
        RECT 526.290000 298.620000 527.090000 299.100000 ;
        RECT 526.290000 304.060000 527.090000 304.540000 ;
        RECT 526.290000 325.820000 527.090000 326.300000 ;
        RECT 526.290000 309.500000 527.090000 309.980000 ;
        RECT 526.290000 314.940000 527.090000 315.420000 ;
        RECT 526.290000 320.380000 527.090000 320.860000 ;
        RECT 526.290000 336.700000 527.090000 337.180000 ;
        RECT 526.290000 331.260000 527.090000 331.740000 ;
        RECT 526.290000 347.580000 527.090000 348.060000 ;
        RECT 526.290000 353.020000 527.090000 353.500000 ;
        RECT 526.290000 358.460000 527.090000 358.940000 ;
        RECT 526.290000 363.900000 527.090000 364.380000 ;
        RECT 526.290000 369.340000 527.090000 369.820000 ;
        RECT 526.290000 374.780000 527.090000 375.260000 ;
        RECT 526.290000 380.220000 527.090000 380.700000 ;
        RECT 526.290000 385.660000 527.090000 386.140000 ;
        RECT 526.290000 391.100000 527.090000 391.580000 ;
        RECT 526.290000 396.540000 527.090000 397.020000 ;
        RECT 526.290000 401.980000 527.090000 402.460000 ;
        RECT 526.290000 407.420000 527.090000 407.900000 ;
        RECT 526.290000 412.860000 527.090000 413.340000 ;
      LAYER met4 ;
        RECT 526.290000 0.000000 527.090000 420.240000 ;
        RECT 2.830000 0.000000 3.630000 420.240000 ;
    END
# end of P/G power stripe data as pin


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 34.820000 403.640000 505.080000 405.380000 ;
      LAYER met3 ;
        RECT 34.820000 17.400000 505.080000 19.140000 ;
      LAYER met4 ;
        RECT 34.820000 17.400000 36.560000 405.380000 ;
      LAYER met4 ;
        RECT 503.340000 17.400000 505.080000 405.380000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 529.120000 416.970000 529.920000 417.770000 ;
    END
    PORT
      LAYER met3 ;
        RECT 529.120000 1.450000 529.920000 2.250000 ;
    END
    PORT
      LAYER met4 ;
        RECT 527.690000 419.440000 528.490000 420.240000 ;
    END
    PORT
      LAYER met4 ;
        RECT 527.690000 0.000000 528.490000 0.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.430000 419.440000 2.230000 420.240000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.430000 0.000000 2.230000 0.800000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 1.430000 1.450000 529.920000 2.250000 ;
        RECT 1.430000 416.970000 529.920000 417.770000 ;
        RECT 1.430000 7.580000 2.230000 8.060000 ;
        RECT 1.430000 13.020000 2.230000 13.500000 ;
        RECT 1.430000 18.460000 2.230000 18.940000 ;
        RECT 1.430000 23.900000 2.230000 24.380000 ;
        RECT 1.430000 29.340000 2.230000 29.820000 ;
        RECT 1.430000 34.780000 2.230000 35.260000 ;
        RECT 1.430000 40.220000 2.230000 40.700000 ;
        RECT 1.430000 45.660000 2.230000 46.140000 ;
        RECT 1.430000 51.100000 2.230000 51.580000 ;
        RECT 1.430000 56.540000 2.230000 57.020000 ;
        RECT 1.430000 61.980000 2.230000 62.460000 ;
        RECT 1.430000 67.420000 2.230000 67.900000 ;
        RECT 1.430000 72.860000 2.230000 73.340000 ;
        RECT 1.430000 143.580000 2.230000 144.060000 ;
        RECT 1.430000 78.300000 2.230000 78.780000 ;
        RECT 1.430000 83.740000 2.230000 84.220000 ;
        RECT 1.430000 89.180000 2.230000 89.660000 ;
        RECT 1.430000 94.620000 2.230000 95.100000 ;
        RECT 1.430000 100.060000 2.230000 100.540000 ;
        RECT 1.430000 105.500000 2.230000 105.980000 ;
        RECT 1.430000 127.260000 2.230000 127.740000 ;
        RECT 1.430000 110.940000 2.230000 111.420000 ;
        RECT 1.430000 116.380000 2.230000 116.860000 ;
        RECT 1.430000 121.820000 2.230000 122.300000 ;
        RECT 1.430000 138.140000 2.230000 138.620000 ;
        RECT 1.430000 132.700000 2.230000 133.180000 ;
        RECT 1.430000 149.020000 2.230000 149.500000 ;
        RECT 1.430000 154.460000 2.230000 154.940000 ;
        RECT 1.430000 159.900000 2.230000 160.380000 ;
        RECT 1.430000 165.340000 2.230000 165.820000 ;
        RECT 1.430000 170.780000 2.230000 171.260000 ;
        RECT 1.430000 176.220000 2.230000 176.700000 ;
        RECT 1.430000 181.660000 2.230000 182.140000 ;
        RECT 1.430000 187.100000 2.230000 187.580000 ;
        RECT 1.430000 192.540000 2.230000 193.020000 ;
        RECT 1.430000 197.980000 2.230000 198.460000 ;
        RECT 1.430000 203.420000 2.230000 203.900000 ;
        RECT 1.430000 208.860000 2.230000 209.340000 ;
        RECT 527.690000 7.580000 528.490000 8.060000 ;
        RECT 527.690000 13.020000 528.490000 13.500000 ;
        RECT 527.690000 18.460000 528.490000 18.940000 ;
        RECT 527.690000 23.900000 528.490000 24.380000 ;
        RECT 527.690000 29.340000 528.490000 29.820000 ;
        RECT 527.690000 34.780000 528.490000 35.260000 ;
        RECT 527.690000 40.220000 528.490000 40.700000 ;
        RECT 527.690000 45.660000 528.490000 46.140000 ;
        RECT 527.690000 51.100000 528.490000 51.580000 ;
        RECT 527.690000 56.540000 528.490000 57.020000 ;
        RECT 527.690000 61.980000 528.490000 62.460000 ;
        RECT 527.690000 67.420000 528.490000 67.900000 ;
        RECT 527.690000 72.860000 528.490000 73.340000 ;
        RECT 527.690000 143.580000 528.490000 144.060000 ;
        RECT 527.690000 78.300000 528.490000 78.780000 ;
        RECT 527.690000 83.740000 528.490000 84.220000 ;
        RECT 527.690000 89.180000 528.490000 89.660000 ;
        RECT 527.690000 94.620000 528.490000 95.100000 ;
        RECT 527.690000 100.060000 528.490000 100.540000 ;
        RECT 527.690000 105.500000 528.490000 105.980000 ;
        RECT 527.690000 127.260000 528.490000 127.740000 ;
        RECT 527.690000 110.940000 528.490000 111.420000 ;
        RECT 527.690000 116.380000 528.490000 116.860000 ;
        RECT 527.690000 121.820000 528.490000 122.300000 ;
        RECT 527.690000 138.140000 528.490000 138.620000 ;
        RECT 527.690000 132.700000 528.490000 133.180000 ;
        RECT 527.690000 149.020000 528.490000 149.500000 ;
        RECT 527.690000 154.460000 528.490000 154.940000 ;
        RECT 527.690000 159.900000 528.490000 160.380000 ;
        RECT 527.690000 165.340000 528.490000 165.820000 ;
        RECT 527.690000 170.780000 528.490000 171.260000 ;
        RECT 527.690000 176.220000 528.490000 176.700000 ;
        RECT 527.690000 181.660000 528.490000 182.140000 ;
        RECT 527.690000 187.100000 528.490000 187.580000 ;
        RECT 527.690000 192.540000 528.490000 193.020000 ;
        RECT 527.690000 197.980000 528.490000 198.460000 ;
        RECT 527.690000 203.420000 528.490000 203.900000 ;
        RECT 527.690000 208.860000 528.490000 209.340000 ;
        RECT 1.430000 214.300000 2.230000 214.780000 ;
        RECT 1.430000 219.740000 2.230000 220.220000 ;
        RECT 1.430000 225.180000 2.230000 225.660000 ;
        RECT 1.430000 230.620000 2.230000 231.100000 ;
        RECT 1.430000 236.060000 2.230000 236.540000 ;
        RECT 1.430000 241.500000 2.230000 241.980000 ;
        RECT 1.430000 246.940000 2.230000 247.420000 ;
        RECT 1.430000 252.380000 2.230000 252.860000 ;
        RECT 1.430000 257.820000 2.230000 258.300000 ;
        RECT 1.430000 263.260000 2.230000 263.740000 ;
        RECT 1.430000 268.700000 2.230000 269.180000 ;
        RECT 1.430000 274.140000 2.230000 274.620000 ;
        RECT 1.430000 279.580000 2.230000 280.060000 ;
        RECT 1.430000 285.020000 2.230000 285.500000 ;
        RECT 1.430000 290.460000 2.230000 290.940000 ;
        RECT 1.430000 295.900000 2.230000 296.380000 ;
        RECT 1.430000 301.340000 2.230000 301.820000 ;
        RECT 1.430000 306.780000 2.230000 307.260000 ;
        RECT 1.430000 312.220000 2.230000 312.700000 ;
        RECT 1.430000 317.660000 2.230000 318.140000 ;
        RECT 1.430000 323.100000 2.230000 323.580000 ;
        RECT 1.430000 339.420000 2.230000 339.900000 ;
        RECT 1.430000 333.980000 2.230000 334.460000 ;
        RECT 1.430000 328.540000 2.230000 329.020000 ;
        RECT 1.430000 344.860000 2.230000 345.340000 ;
        RECT 1.430000 350.300000 2.230000 350.780000 ;
        RECT 1.430000 355.740000 2.230000 356.220000 ;
        RECT 1.430000 361.180000 2.230000 361.660000 ;
        RECT 1.430000 366.620000 2.230000 367.100000 ;
        RECT 1.430000 372.060000 2.230000 372.540000 ;
        RECT 1.430000 377.500000 2.230000 377.980000 ;
        RECT 1.430000 382.940000 2.230000 383.420000 ;
        RECT 1.430000 388.380000 2.230000 388.860000 ;
        RECT 1.430000 393.820000 2.230000 394.300000 ;
        RECT 1.430000 399.260000 2.230000 399.740000 ;
        RECT 1.430000 404.700000 2.230000 405.180000 ;
        RECT 1.430000 410.140000 2.230000 410.620000 ;
        RECT 527.690000 214.300000 528.490000 214.780000 ;
        RECT 527.690000 219.740000 528.490000 220.220000 ;
        RECT 527.690000 225.180000 528.490000 225.660000 ;
        RECT 527.690000 230.620000 528.490000 231.100000 ;
        RECT 527.690000 236.060000 528.490000 236.540000 ;
        RECT 527.690000 241.500000 528.490000 241.980000 ;
        RECT 527.690000 246.940000 528.490000 247.420000 ;
        RECT 527.690000 252.380000 528.490000 252.860000 ;
        RECT 527.690000 257.820000 528.490000 258.300000 ;
        RECT 527.690000 263.260000 528.490000 263.740000 ;
        RECT 527.690000 268.700000 528.490000 269.180000 ;
        RECT 527.690000 274.140000 528.490000 274.620000 ;
        RECT 527.690000 279.580000 528.490000 280.060000 ;
        RECT 527.690000 285.020000 528.490000 285.500000 ;
        RECT 527.690000 290.460000 528.490000 290.940000 ;
        RECT 527.690000 295.900000 528.490000 296.380000 ;
        RECT 527.690000 301.340000 528.490000 301.820000 ;
        RECT 527.690000 306.780000 528.490000 307.260000 ;
        RECT 527.690000 312.220000 528.490000 312.700000 ;
        RECT 527.690000 317.660000 528.490000 318.140000 ;
        RECT 527.690000 323.100000 528.490000 323.580000 ;
        RECT 527.690000 339.420000 528.490000 339.900000 ;
        RECT 527.690000 333.980000 528.490000 334.460000 ;
        RECT 527.690000 328.540000 528.490000 329.020000 ;
        RECT 527.690000 344.860000 528.490000 345.340000 ;
        RECT 527.690000 350.300000 528.490000 350.780000 ;
        RECT 527.690000 355.740000 528.490000 356.220000 ;
        RECT 527.690000 361.180000 528.490000 361.660000 ;
        RECT 527.690000 366.620000 528.490000 367.100000 ;
        RECT 527.690000 372.060000 528.490000 372.540000 ;
        RECT 527.690000 377.500000 528.490000 377.980000 ;
        RECT 527.690000 382.940000 528.490000 383.420000 ;
        RECT 527.690000 388.380000 528.490000 388.860000 ;
        RECT 527.690000 393.820000 528.490000 394.300000 ;
        RECT 527.690000 399.260000 528.490000 399.740000 ;
        RECT 527.690000 404.700000 528.490000 405.180000 ;
        RECT 527.690000 410.140000 528.490000 410.620000 ;
      LAYER met4 ;
        RECT 527.690000 0.000000 528.490000 420.240000 ;
        RECT 1.430000 0.000000 2.230000 420.240000 ;
    END
# end of P/G power stripe data as pin


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 506.740000 14.000000 508.480000 408.780000 ;
      LAYER met3 ;
        RECT 31.420000 14.000000 508.480000 15.740000 ;
      LAYER met3 ;
        RECT 31.420000 407.040000 508.480000 408.780000 ;
      LAYER met4 ;
        RECT 31.420000 14.000000 33.160000 408.780000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 529.920000 420.240000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 529.920000 420.240000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 529.920000 420.240000 ;
    LAYER met3 ;
      RECT 0.000000 418.070000 529.920000 420.240000 ;
      RECT 0.000000 416.670000 1.130000 418.070000 ;
      RECT 0.000000 415.270000 2.530000 416.670000 ;
      RECT 0.000000 413.640000 529.920000 415.270000 ;
      RECT 527.390000 412.560000 529.920000 413.640000 ;
      RECT 3.930000 412.560000 525.990000 413.640000 ;
      RECT 0.000000 412.560000 2.530000 413.640000 ;
      RECT 0.000000 410.920000 529.920000 412.560000 ;
      RECT 528.790000 409.840000 529.920000 410.920000 ;
      RECT 2.530000 409.840000 527.390000 410.920000 ;
      RECT 0.000000 409.840000 1.130000 410.920000 ;
      RECT 0.000000 408.200000 529.920000 409.840000 ;
      RECT 527.390000 407.120000 529.920000 408.200000 ;
      RECT 3.930000 407.120000 525.990000 408.200000 ;
      RECT 0.000000 407.120000 2.530000 408.200000 ;
      RECT 0.000000 405.480000 529.920000 407.120000 ;
      RECT 528.790000 404.400000 529.920000 405.480000 ;
      RECT 2.530000 404.400000 527.390000 405.480000 ;
      RECT 0.000000 404.400000 1.130000 405.480000 ;
      RECT 0.000000 402.760000 529.920000 404.400000 ;
      RECT 527.390000 401.680000 529.920000 402.760000 ;
      RECT 3.930000 401.680000 525.990000 402.760000 ;
      RECT 0.000000 401.680000 2.530000 402.760000 ;
      RECT 0.000000 400.040000 529.920000 401.680000 ;
      RECT 0.000000 399.820000 1.130000 400.040000 ;
      RECT 528.790000 398.960000 529.920000 400.040000 ;
      RECT 2.530000 398.960000 527.390000 400.040000 ;
      RECT 1.020000 398.960000 1.130000 399.820000 ;
      RECT 1.020000 398.840000 529.920000 398.960000 ;
      RECT 0.000000 397.320000 529.920000 398.840000 ;
      RECT 527.390000 396.240000 529.920000 397.320000 ;
      RECT 3.930000 396.240000 525.990000 397.320000 ;
      RECT 0.000000 396.240000 2.530000 397.320000 ;
      RECT 0.000000 395.550000 529.920000 396.240000 ;
      RECT 1.020000 394.600000 529.920000 395.550000 ;
      RECT 1.020000 394.570000 1.130000 394.600000 ;
      RECT 528.790000 393.520000 529.920000 394.600000 ;
      RECT 2.530000 393.520000 527.390000 394.600000 ;
      RECT 0.000000 393.520000 1.130000 394.570000 ;
      RECT 0.000000 391.880000 529.920000 393.520000 ;
      RECT 527.390000 390.800000 529.920000 391.880000 ;
      RECT 3.930000 390.800000 525.990000 391.880000 ;
      RECT 0.000000 390.800000 2.530000 391.880000 ;
      RECT 0.000000 390.670000 529.920000 390.800000 ;
      RECT 1.020000 389.690000 529.920000 390.670000 ;
      RECT 0.000000 389.160000 529.920000 389.690000 ;
      RECT 528.790000 388.080000 529.920000 389.160000 ;
      RECT 2.530000 388.080000 527.390000 389.160000 ;
      RECT 0.000000 388.080000 1.130000 389.160000 ;
      RECT 0.000000 386.440000 529.920000 388.080000 ;
      RECT 0.000000 385.790000 2.530000 386.440000 ;
      RECT 527.390000 385.360000 529.920000 386.440000 ;
      RECT 3.930000 385.360000 525.990000 386.440000 ;
      RECT 1.020000 385.360000 2.530000 385.790000 ;
      RECT 1.020000 384.810000 529.920000 385.360000 ;
      RECT 0.000000 383.720000 529.920000 384.810000 ;
      RECT 528.790000 382.640000 529.920000 383.720000 ;
      RECT 2.530000 382.640000 527.390000 383.720000 ;
      RECT 0.000000 382.640000 1.130000 383.720000 ;
      RECT 0.000000 381.000000 529.920000 382.640000 ;
      RECT 0.000000 380.910000 2.530000 381.000000 ;
      RECT 1.020000 379.930000 2.530000 380.910000 ;
      RECT 527.390000 379.920000 529.920000 381.000000 ;
      RECT 3.930000 379.920000 525.990000 381.000000 ;
      RECT 0.000000 379.920000 2.530000 379.930000 ;
      RECT 0.000000 378.280000 529.920000 379.920000 ;
      RECT 528.790000 377.200000 529.920000 378.280000 ;
      RECT 2.530000 377.200000 527.390000 378.280000 ;
      RECT 0.000000 377.200000 1.130000 378.280000 ;
      RECT 0.000000 376.640000 529.920000 377.200000 ;
      RECT 1.020000 375.660000 529.920000 376.640000 ;
      RECT 0.000000 375.560000 529.920000 375.660000 ;
      RECT 527.390000 374.480000 529.920000 375.560000 ;
      RECT 3.930000 374.480000 525.990000 375.560000 ;
      RECT 0.000000 374.480000 2.530000 375.560000 ;
      RECT 0.000000 372.840000 529.920000 374.480000 ;
      RECT 528.790000 371.760000 529.920000 372.840000 ;
      RECT 2.530000 371.760000 527.390000 372.840000 ;
      RECT 0.000000 371.760000 1.130000 372.840000 ;
      RECT 1.020000 370.780000 529.920000 371.760000 ;
      RECT 0.000000 370.120000 529.920000 370.780000 ;
      RECT 527.390000 369.040000 529.920000 370.120000 ;
      RECT 3.930000 369.040000 525.990000 370.120000 ;
      RECT 0.000000 369.040000 2.530000 370.120000 ;
      RECT 0.000000 367.400000 529.920000 369.040000 ;
      RECT 0.000000 366.880000 1.130000 367.400000 ;
      RECT 528.790000 366.320000 529.920000 367.400000 ;
      RECT 2.530000 366.320000 527.390000 367.400000 ;
      RECT 1.020000 366.320000 1.130000 366.880000 ;
      RECT 1.020000 365.900000 529.920000 366.320000 ;
      RECT 0.000000 364.680000 529.920000 365.900000 ;
      RECT 527.390000 363.600000 529.920000 364.680000 ;
      RECT 3.930000 363.600000 525.990000 364.680000 ;
      RECT 0.000000 363.600000 2.530000 364.680000 ;
      RECT 0.000000 362.000000 529.920000 363.600000 ;
      RECT 1.020000 361.960000 529.920000 362.000000 ;
      RECT 1.020000 361.020000 1.130000 361.960000 ;
      RECT 528.790000 360.880000 529.920000 361.960000 ;
      RECT 2.530000 360.880000 527.390000 361.960000 ;
      RECT 0.000000 360.880000 1.130000 361.020000 ;
      RECT 0.000000 359.240000 529.920000 360.880000 ;
      RECT 527.390000 358.160000 529.920000 359.240000 ;
      RECT 3.930000 358.160000 525.990000 359.240000 ;
      RECT 0.000000 358.160000 2.530000 359.240000 ;
      RECT 0.000000 357.120000 529.920000 358.160000 ;
      RECT 1.020000 356.520000 529.920000 357.120000 ;
      RECT 1.020000 356.140000 1.130000 356.520000 ;
      RECT 528.790000 355.440000 529.920000 356.520000 ;
      RECT 2.530000 355.440000 527.390000 356.520000 ;
      RECT 0.000000 355.440000 1.130000 356.140000 ;
      RECT 0.000000 353.800000 529.920000 355.440000 ;
      RECT 0.000000 352.850000 2.530000 353.800000 ;
      RECT 527.390000 352.720000 529.920000 353.800000 ;
      RECT 3.930000 352.720000 525.990000 353.800000 ;
      RECT 1.020000 352.720000 2.530000 352.850000 ;
      RECT 1.020000 351.870000 529.920000 352.720000 ;
      RECT 0.000000 351.080000 529.920000 351.870000 ;
      RECT 528.790000 350.000000 529.920000 351.080000 ;
      RECT 2.530000 350.000000 527.390000 351.080000 ;
      RECT 0.000000 350.000000 1.130000 351.080000 ;
      RECT 0.000000 348.360000 529.920000 350.000000 ;
      RECT 0.000000 347.970000 2.530000 348.360000 ;
      RECT 527.390000 347.280000 529.920000 348.360000 ;
      RECT 3.930000 347.280000 525.990000 348.360000 ;
      RECT 1.020000 347.280000 2.530000 347.970000 ;
      RECT 1.020000 346.990000 529.920000 347.280000 ;
      RECT 0.000000 345.640000 529.920000 346.990000 ;
      RECT 528.790000 344.560000 529.920000 345.640000 ;
      RECT 2.530000 344.560000 527.390000 345.640000 ;
      RECT 0.000000 344.560000 1.130000 345.640000 ;
      RECT 0.000000 343.090000 529.920000 344.560000 ;
      RECT 1.020000 342.920000 529.920000 343.090000 ;
      RECT 1.020000 342.110000 2.530000 342.920000 ;
      RECT 527.390000 341.840000 529.920000 342.920000 ;
      RECT 3.930000 341.840000 525.990000 342.920000 ;
      RECT 0.000000 341.840000 2.530000 342.110000 ;
      RECT 0.000000 340.200000 529.920000 341.840000 ;
      RECT 528.790000 339.120000 529.920000 340.200000 ;
      RECT 2.530000 339.120000 527.390000 340.200000 ;
      RECT 0.000000 339.120000 1.130000 340.200000 ;
      RECT 0.000000 338.210000 529.920000 339.120000 ;
      RECT 1.020000 337.480000 529.920000 338.210000 ;
      RECT 1.020000 337.230000 2.530000 337.480000 ;
      RECT 527.390000 336.400000 529.920000 337.480000 ;
      RECT 3.930000 336.400000 525.990000 337.480000 ;
      RECT 0.000000 336.400000 2.530000 337.230000 ;
      RECT 0.000000 334.760000 529.920000 336.400000 ;
      RECT 0.000000 333.940000 1.130000 334.760000 ;
      RECT 528.790000 333.680000 529.920000 334.760000 ;
      RECT 2.530000 333.680000 527.390000 334.760000 ;
      RECT 1.020000 333.680000 1.130000 333.940000 ;
      RECT 1.020000 332.960000 529.920000 333.680000 ;
      RECT 0.000000 332.040000 529.920000 332.960000 ;
      RECT 527.390000 330.960000 529.920000 332.040000 ;
      RECT 3.930000 330.960000 525.990000 332.040000 ;
      RECT 0.000000 330.960000 2.530000 332.040000 ;
      RECT 0.000000 329.320000 529.920000 330.960000 ;
      RECT 0.000000 329.060000 1.130000 329.320000 ;
      RECT 528.790000 328.240000 529.920000 329.320000 ;
      RECT 2.530000 328.240000 527.390000 329.320000 ;
      RECT 1.020000 328.240000 1.130000 329.060000 ;
      RECT 1.020000 328.080000 529.920000 328.240000 ;
      RECT 0.000000 326.600000 529.920000 328.080000 ;
      RECT 527.390000 325.520000 529.920000 326.600000 ;
      RECT 3.930000 325.520000 525.990000 326.600000 ;
      RECT 0.000000 325.520000 2.530000 326.600000 ;
      RECT 0.000000 324.180000 529.920000 325.520000 ;
      RECT 1.020000 323.880000 529.920000 324.180000 ;
      RECT 1.020000 323.200000 1.130000 323.880000 ;
      RECT 528.790000 322.800000 529.920000 323.880000 ;
      RECT 2.530000 322.800000 527.390000 323.880000 ;
      RECT 0.000000 322.800000 1.130000 323.200000 ;
      RECT 0.000000 321.160000 529.920000 322.800000 ;
      RECT 527.390000 320.080000 529.920000 321.160000 ;
      RECT 3.930000 320.080000 525.990000 321.160000 ;
      RECT 0.000000 320.080000 2.530000 321.160000 ;
      RECT 0.000000 319.300000 529.920000 320.080000 ;
      RECT 1.020000 318.440000 529.920000 319.300000 ;
      RECT 1.020000 318.320000 1.130000 318.440000 ;
      RECT 528.790000 317.360000 529.920000 318.440000 ;
      RECT 2.530000 317.360000 527.390000 318.440000 ;
      RECT 0.000000 317.360000 1.130000 318.320000 ;
      RECT 0.000000 315.720000 529.920000 317.360000 ;
      RECT 527.390000 314.640000 529.920000 315.720000 ;
      RECT 3.930000 314.640000 525.990000 315.720000 ;
      RECT 0.000000 314.640000 2.530000 315.720000 ;
      RECT 0.000000 314.420000 529.920000 314.640000 ;
      RECT 1.020000 313.440000 529.920000 314.420000 ;
      RECT 0.000000 313.000000 529.920000 313.440000 ;
      RECT 528.790000 311.920000 529.920000 313.000000 ;
      RECT 2.530000 311.920000 527.390000 313.000000 ;
      RECT 0.000000 311.920000 1.130000 313.000000 ;
      RECT 0.000000 310.280000 529.920000 311.920000 ;
      RECT 0.000000 310.150000 2.530000 310.280000 ;
      RECT 527.390000 309.200000 529.920000 310.280000 ;
      RECT 3.930000 309.200000 525.990000 310.280000 ;
      RECT 1.020000 309.200000 2.530000 310.150000 ;
      RECT 1.020000 309.170000 529.920000 309.200000 ;
      RECT 0.000000 307.560000 529.920000 309.170000 ;
      RECT 528.790000 306.480000 529.920000 307.560000 ;
      RECT 2.530000 306.480000 527.390000 307.560000 ;
      RECT 0.000000 306.480000 1.130000 307.560000 ;
      RECT 0.000000 305.270000 529.920000 306.480000 ;
      RECT 1.020000 304.840000 529.920000 305.270000 ;
      RECT 1.020000 304.290000 2.530000 304.840000 ;
      RECT 527.390000 303.760000 529.920000 304.840000 ;
      RECT 3.930000 303.760000 525.990000 304.840000 ;
      RECT 0.000000 303.760000 2.530000 304.290000 ;
      RECT 0.000000 302.120000 529.920000 303.760000 ;
      RECT 528.790000 301.040000 529.920000 302.120000 ;
      RECT 2.530000 301.040000 527.390000 302.120000 ;
      RECT 0.000000 301.040000 1.130000 302.120000 ;
      RECT 0.000000 300.390000 529.920000 301.040000 ;
      RECT 1.020000 299.410000 529.920000 300.390000 ;
      RECT 0.000000 299.400000 529.920000 299.410000 ;
      RECT 527.390000 298.320000 529.920000 299.400000 ;
      RECT 3.930000 298.320000 525.990000 299.400000 ;
      RECT 0.000000 298.320000 2.530000 299.400000 ;
      RECT 0.000000 296.680000 529.920000 298.320000 ;
      RECT 528.790000 295.600000 529.920000 296.680000 ;
      RECT 2.530000 295.600000 527.390000 296.680000 ;
      RECT 0.000000 295.600000 1.130000 296.680000 ;
      RECT 0.000000 295.510000 529.920000 295.600000 ;
      RECT 1.020000 294.530000 529.920000 295.510000 ;
      RECT 0.000000 293.960000 529.920000 294.530000 ;
      RECT 527.390000 292.880000 529.920000 293.960000 ;
      RECT 3.930000 292.880000 525.990000 293.960000 ;
      RECT 0.000000 292.880000 2.530000 293.960000 ;
      RECT 0.000000 291.240000 529.920000 292.880000 ;
      RECT 1.020000 290.260000 1.130000 291.240000 ;
      RECT 528.790000 290.160000 529.920000 291.240000 ;
      RECT 2.530000 290.160000 527.390000 291.240000 ;
      RECT 0.000000 290.160000 1.130000 290.260000 ;
      RECT 0.000000 288.520000 529.920000 290.160000 ;
      RECT 527.390000 287.440000 529.920000 288.520000 ;
      RECT 3.930000 287.440000 525.990000 288.520000 ;
      RECT 0.000000 287.440000 2.530000 288.520000 ;
      RECT 0.000000 286.360000 529.920000 287.440000 ;
      RECT 1.020000 285.800000 529.920000 286.360000 ;
      RECT 1.020000 285.380000 1.130000 285.800000 ;
      RECT 528.790000 284.720000 529.920000 285.800000 ;
      RECT 2.530000 284.720000 527.390000 285.800000 ;
      RECT 0.000000 284.720000 1.130000 285.380000 ;
      RECT 0.000000 283.080000 529.920000 284.720000 ;
      RECT 527.390000 282.000000 529.920000 283.080000 ;
      RECT 3.930000 282.000000 525.990000 283.080000 ;
      RECT 0.000000 282.000000 2.530000 283.080000 ;
      RECT 0.000000 281.480000 529.920000 282.000000 ;
      RECT 1.020000 280.500000 529.920000 281.480000 ;
      RECT 0.000000 280.360000 529.920000 280.500000 ;
      RECT 528.790000 279.280000 529.920000 280.360000 ;
      RECT 2.530000 279.280000 527.390000 280.360000 ;
      RECT 0.000000 279.280000 1.130000 280.360000 ;
      RECT 0.000000 277.640000 529.920000 279.280000 ;
      RECT 0.000000 276.600000 2.530000 277.640000 ;
      RECT 527.390000 276.560000 529.920000 277.640000 ;
      RECT 3.930000 276.560000 525.990000 277.640000 ;
      RECT 1.020000 276.560000 2.530000 276.600000 ;
      RECT 1.020000 275.620000 529.920000 276.560000 ;
      RECT 0.000000 274.920000 529.920000 275.620000 ;
      RECT 528.790000 273.840000 529.920000 274.920000 ;
      RECT 2.530000 273.840000 527.390000 274.920000 ;
      RECT 0.000000 273.840000 1.130000 274.920000 ;
      RECT 0.000000 272.200000 529.920000 273.840000 ;
      RECT 0.000000 271.720000 2.530000 272.200000 ;
      RECT 527.390000 271.120000 529.920000 272.200000 ;
      RECT 3.930000 271.120000 525.990000 272.200000 ;
      RECT 1.020000 271.120000 2.530000 271.720000 ;
      RECT 1.020000 270.740000 529.920000 271.120000 ;
      RECT 0.000000 269.480000 529.920000 270.740000 ;
      RECT 528.790000 268.400000 529.920000 269.480000 ;
      RECT 2.530000 268.400000 527.390000 269.480000 ;
      RECT 0.000000 268.400000 1.130000 269.480000 ;
      RECT 0.000000 267.450000 529.920000 268.400000 ;
      RECT 1.020000 266.760000 529.920000 267.450000 ;
      RECT 1.020000 266.470000 2.530000 266.760000 ;
      RECT 527.390000 265.680000 529.920000 266.760000 ;
      RECT 3.930000 265.680000 525.990000 266.760000 ;
      RECT 0.000000 265.680000 2.530000 266.470000 ;
      RECT 0.000000 264.040000 529.920000 265.680000 ;
      RECT 528.790000 262.960000 529.920000 264.040000 ;
      RECT 2.530000 262.960000 527.390000 264.040000 ;
      RECT 0.000000 262.960000 1.130000 264.040000 ;
      RECT 0.000000 262.570000 529.920000 262.960000 ;
      RECT 1.020000 261.590000 529.920000 262.570000 ;
      RECT 0.000000 261.320000 529.920000 261.590000 ;
      RECT 527.390000 260.240000 529.920000 261.320000 ;
      RECT 3.930000 260.240000 525.990000 261.320000 ;
      RECT 0.000000 260.240000 2.530000 261.320000 ;
      RECT 0.000000 258.600000 529.920000 260.240000 ;
      RECT 0.000000 257.690000 1.130000 258.600000 ;
      RECT 528.790000 257.520000 529.920000 258.600000 ;
      RECT 2.530000 257.520000 527.390000 258.600000 ;
      RECT 1.020000 257.520000 1.130000 257.690000 ;
      RECT 1.020000 256.710000 529.920000 257.520000 ;
      RECT 0.000000 255.880000 529.920000 256.710000 ;
      RECT 527.390000 254.800000 529.920000 255.880000 ;
      RECT 3.930000 254.800000 525.990000 255.880000 ;
      RECT 0.000000 254.800000 2.530000 255.880000 ;
      RECT 0.000000 253.160000 529.920000 254.800000 ;
      RECT 0.000000 252.810000 1.130000 253.160000 ;
      RECT 528.790000 252.080000 529.920000 253.160000 ;
      RECT 2.530000 252.080000 527.390000 253.160000 ;
      RECT 1.020000 252.080000 1.130000 252.810000 ;
      RECT 1.020000 251.830000 529.920000 252.080000 ;
      RECT 0.000000 250.440000 529.920000 251.830000 ;
      RECT 527.390000 249.360000 529.920000 250.440000 ;
      RECT 3.930000 249.360000 525.990000 250.440000 ;
      RECT 0.000000 249.360000 2.530000 250.440000 ;
      RECT 0.000000 248.540000 529.920000 249.360000 ;
      RECT 1.020000 247.720000 529.920000 248.540000 ;
      RECT 1.020000 247.560000 1.130000 247.720000 ;
      RECT 528.790000 246.640000 529.920000 247.720000 ;
      RECT 2.530000 246.640000 527.390000 247.720000 ;
      RECT 0.000000 246.640000 1.130000 247.560000 ;
      RECT 0.000000 245.000000 529.920000 246.640000 ;
      RECT 527.390000 243.920000 529.920000 245.000000 ;
      RECT 3.930000 243.920000 525.990000 245.000000 ;
      RECT 0.000000 243.920000 2.530000 245.000000 ;
      RECT 0.000000 243.660000 529.920000 243.920000 ;
      RECT 1.020000 242.680000 529.920000 243.660000 ;
      RECT 0.000000 242.280000 529.920000 242.680000 ;
      RECT 528.790000 241.200000 529.920000 242.280000 ;
      RECT 2.530000 241.200000 527.390000 242.280000 ;
      RECT 0.000000 241.200000 1.130000 242.280000 ;
      RECT 0.000000 239.560000 529.920000 241.200000 ;
      RECT 0.000000 238.780000 2.530000 239.560000 ;
      RECT 527.390000 238.480000 529.920000 239.560000 ;
      RECT 3.930000 238.480000 525.990000 239.560000 ;
      RECT 1.020000 238.480000 2.530000 238.780000 ;
      RECT 1.020000 237.800000 529.920000 238.480000 ;
      RECT 0.000000 236.840000 529.920000 237.800000 ;
      RECT 528.790000 235.760000 529.920000 236.840000 ;
      RECT 2.530000 235.760000 527.390000 236.840000 ;
      RECT 0.000000 235.760000 1.130000 236.840000 ;
      RECT 0.000000 234.120000 529.920000 235.760000 ;
      RECT 0.000000 233.900000 2.530000 234.120000 ;
      RECT 527.390000 233.040000 529.920000 234.120000 ;
      RECT 3.930000 233.040000 525.990000 234.120000 ;
      RECT 1.020000 233.040000 2.530000 233.900000 ;
      RECT 1.020000 232.920000 529.920000 233.040000 ;
      RECT 0.000000 231.400000 529.920000 232.920000 ;
      RECT 528.790000 230.320000 529.920000 231.400000 ;
      RECT 2.530000 230.320000 527.390000 231.400000 ;
      RECT 0.000000 230.320000 1.130000 231.400000 ;
      RECT 0.000000 229.020000 529.920000 230.320000 ;
      RECT 1.020000 228.680000 529.920000 229.020000 ;
      RECT 1.020000 228.040000 2.530000 228.680000 ;
      RECT 527.390000 227.600000 529.920000 228.680000 ;
      RECT 3.930000 227.600000 525.990000 228.680000 ;
      RECT 0.000000 227.600000 2.530000 228.040000 ;
      RECT 0.000000 225.960000 529.920000 227.600000 ;
      RECT 528.790000 224.880000 529.920000 225.960000 ;
      RECT 2.530000 224.880000 527.390000 225.960000 ;
      RECT 0.000000 224.880000 1.130000 225.960000 ;
      RECT 0.000000 224.750000 529.920000 224.880000 ;
      RECT 1.020000 223.770000 529.920000 224.750000 ;
      RECT 0.000000 223.240000 529.920000 223.770000 ;
      RECT 527.390000 222.160000 529.920000 223.240000 ;
      RECT 3.930000 222.160000 525.990000 223.240000 ;
      RECT 0.000000 222.160000 2.530000 223.240000 ;
      RECT 0.000000 220.520000 529.920000 222.160000 ;
      RECT 0.000000 219.870000 1.130000 220.520000 ;
      RECT 528.790000 219.440000 529.920000 220.520000 ;
      RECT 2.530000 219.440000 527.390000 220.520000 ;
      RECT 1.020000 219.440000 1.130000 219.870000 ;
      RECT 1.020000 218.890000 529.920000 219.440000 ;
      RECT 0.000000 217.800000 529.920000 218.890000 ;
      RECT 527.390000 216.720000 529.920000 217.800000 ;
      RECT 3.930000 216.720000 525.990000 217.800000 ;
      RECT 0.000000 216.720000 2.530000 217.800000 ;
      RECT 0.000000 215.080000 529.920000 216.720000 ;
      RECT 0.000000 214.990000 1.130000 215.080000 ;
      RECT 1.020000 214.010000 1.130000 214.990000 ;
      RECT 528.790000 214.000000 529.920000 215.080000 ;
      RECT 2.530000 214.000000 527.390000 215.080000 ;
      RECT 0.000000 214.000000 1.130000 214.010000 ;
      RECT 0.000000 212.360000 529.920000 214.000000 ;
      RECT 527.390000 211.280000 529.920000 212.360000 ;
      RECT 3.930000 211.280000 525.990000 212.360000 ;
      RECT 0.000000 211.280000 2.530000 212.360000 ;
      RECT 0.000000 210.110000 529.920000 211.280000 ;
      RECT 1.020000 209.640000 529.920000 210.110000 ;
      RECT 1.020000 209.130000 1.130000 209.640000 ;
      RECT 528.790000 208.560000 529.920000 209.640000 ;
      RECT 2.530000 208.560000 527.390000 209.640000 ;
      RECT 0.000000 208.560000 1.130000 209.130000 ;
      RECT 0.000000 206.920000 529.920000 208.560000 ;
      RECT 527.390000 205.840000 529.920000 206.920000 ;
      RECT 3.930000 205.840000 525.990000 206.920000 ;
      RECT 0.000000 205.840000 2.530000 206.920000 ;
      RECT 1.020000 204.860000 529.920000 205.840000 ;
      RECT 0.000000 204.200000 529.920000 204.860000 ;
      RECT 528.790000 203.120000 529.920000 204.200000 ;
      RECT 2.530000 203.120000 527.390000 204.200000 ;
      RECT 0.000000 203.120000 1.130000 204.200000 ;
      RECT 0.000000 201.480000 529.920000 203.120000 ;
      RECT 0.000000 200.960000 2.530000 201.480000 ;
      RECT 527.390000 200.400000 529.920000 201.480000 ;
      RECT 3.930000 200.400000 525.990000 201.480000 ;
      RECT 1.020000 200.400000 2.530000 200.960000 ;
      RECT 1.020000 199.980000 529.920000 200.400000 ;
      RECT 0.000000 198.760000 529.920000 199.980000 ;
      RECT 528.790000 197.680000 529.920000 198.760000 ;
      RECT 2.530000 197.680000 527.390000 198.760000 ;
      RECT 0.000000 197.680000 1.130000 198.760000 ;
      RECT 0.000000 196.040000 529.920000 197.680000 ;
      RECT 527.390000 194.960000 529.920000 196.040000 ;
      RECT 3.930000 194.960000 525.990000 196.040000 ;
      RECT 0.000000 194.960000 2.530000 196.040000 ;
      RECT 0.000000 193.320000 529.920000 194.960000 ;
      RECT 528.790000 192.240000 529.920000 193.320000 ;
      RECT 2.530000 192.240000 527.390000 193.320000 ;
      RECT 0.000000 192.240000 1.130000 193.320000 ;
      RECT 0.000000 190.600000 529.920000 192.240000 ;
      RECT 527.390000 189.520000 529.920000 190.600000 ;
      RECT 3.930000 189.520000 525.990000 190.600000 ;
      RECT 0.000000 189.520000 2.530000 190.600000 ;
      RECT 0.000000 187.880000 529.920000 189.520000 ;
      RECT 528.790000 186.800000 529.920000 187.880000 ;
      RECT 2.530000 186.800000 527.390000 187.880000 ;
      RECT 0.000000 186.800000 1.130000 187.880000 ;
      RECT 0.000000 185.160000 529.920000 186.800000 ;
      RECT 527.390000 184.080000 529.920000 185.160000 ;
      RECT 3.930000 184.080000 525.990000 185.160000 ;
      RECT 0.000000 184.080000 2.530000 185.160000 ;
      RECT 0.000000 182.440000 529.920000 184.080000 ;
      RECT 528.790000 181.360000 529.920000 182.440000 ;
      RECT 2.530000 181.360000 527.390000 182.440000 ;
      RECT 0.000000 181.360000 1.130000 182.440000 ;
      RECT 0.000000 179.720000 529.920000 181.360000 ;
      RECT 527.390000 178.640000 529.920000 179.720000 ;
      RECT 3.930000 178.640000 525.990000 179.720000 ;
      RECT 0.000000 178.640000 2.530000 179.720000 ;
      RECT 0.000000 177.000000 529.920000 178.640000 ;
      RECT 528.790000 175.920000 529.920000 177.000000 ;
      RECT 2.530000 175.920000 527.390000 177.000000 ;
      RECT 0.000000 175.920000 1.130000 177.000000 ;
      RECT 0.000000 174.280000 529.920000 175.920000 ;
      RECT 527.390000 173.200000 529.920000 174.280000 ;
      RECT 3.930000 173.200000 525.990000 174.280000 ;
      RECT 0.000000 173.200000 2.530000 174.280000 ;
      RECT 0.000000 171.560000 529.920000 173.200000 ;
      RECT 528.790000 170.480000 529.920000 171.560000 ;
      RECT 2.530000 170.480000 527.390000 171.560000 ;
      RECT 0.000000 170.480000 1.130000 171.560000 ;
      RECT 0.000000 168.840000 529.920000 170.480000 ;
      RECT 527.390000 167.760000 529.920000 168.840000 ;
      RECT 3.930000 167.760000 525.990000 168.840000 ;
      RECT 0.000000 167.760000 2.530000 168.840000 ;
      RECT 0.000000 166.120000 529.920000 167.760000 ;
      RECT 528.790000 165.040000 529.920000 166.120000 ;
      RECT 2.530000 165.040000 527.390000 166.120000 ;
      RECT 0.000000 165.040000 1.130000 166.120000 ;
      RECT 0.000000 163.400000 529.920000 165.040000 ;
      RECT 527.390000 162.320000 529.920000 163.400000 ;
      RECT 3.930000 162.320000 525.990000 163.400000 ;
      RECT 0.000000 162.320000 2.530000 163.400000 ;
      RECT 0.000000 160.680000 529.920000 162.320000 ;
      RECT 528.790000 159.600000 529.920000 160.680000 ;
      RECT 2.530000 159.600000 527.390000 160.680000 ;
      RECT 0.000000 159.600000 1.130000 160.680000 ;
      RECT 0.000000 157.960000 529.920000 159.600000 ;
      RECT 527.390000 156.880000 529.920000 157.960000 ;
      RECT 3.930000 156.880000 525.990000 157.960000 ;
      RECT 0.000000 156.880000 2.530000 157.960000 ;
      RECT 0.000000 155.240000 529.920000 156.880000 ;
      RECT 528.790000 154.160000 529.920000 155.240000 ;
      RECT 2.530000 154.160000 527.390000 155.240000 ;
      RECT 0.000000 154.160000 1.130000 155.240000 ;
      RECT 0.000000 152.520000 529.920000 154.160000 ;
      RECT 527.390000 151.440000 529.920000 152.520000 ;
      RECT 3.930000 151.440000 525.990000 152.520000 ;
      RECT 0.000000 151.440000 2.530000 152.520000 ;
      RECT 0.000000 149.800000 529.920000 151.440000 ;
      RECT 0.000000 149.720000 1.130000 149.800000 ;
      RECT 1.020000 148.740000 1.130000 149.720000 ;
      RECT 528.790000 148.720000 529.920000 149.800000 ;
      RECT 2.530000 148.720000 527.390000 149.800000 ;
      RECT 0.000000 148.720000 1.130000 148.740000 ;
      RECT 0.000000 147.080000 529.920000 148.720000 ;
      RECT 0.000000 146.670000 2.530000 147.080000 ;
      RECT 527.390000 146.000000 529.920000 147.080000 ;
      RECT 3.930000 146.000000 525.990000 147.080000 ;
      RECT 1.020000 146.000000 2.530000 146.670000 ;
      RECT 1.020000 145.690000 529.920000 146.000000 ;
      RECT 0.000000 144.360000 529.920000 145.690000 ;
      RECT 528.790000 143.280000 529.920000 144.360000 ;
      RECT 2.530000 143.280000 527.390000 144.360000 ;
      RECT 0.000000 143.280000 1.130000 144.360000 ;
      RECT 0.000000 143.010000 529.920000 143.280000 ;
      RECT 1.020000 142.030000 529.920000 143.010000 ;
      RECT 0.000000 141.640000 529.920000 142.030000 ;
      RECT 527.390000 140.560000 529.920000 141.640000 ;
      RECT 3.930000 140.560000 525.990000 141.640000 ;
      RECT 0.000000 140.560000 2.530000 141.640000 ;
      RECT 0.000000 139.960000 529.920000 140.560000 ;
      RECT 1.020000 138.980000 529.920000 139.960000 ;
      RECT 0.000000 138.920000 529.920000 138.980000 ;
      RECT 528.790000 137.840000 529.920000 138.920000 ;
      RECT 2.530000 137.840000 527.390000 138.920000 ;
      RECT 0.000000 137.840000 1.130000 138.920000 ;
      RECT 0.000000 136.300000 529.920000 137.840000 ;
      RECT 1.020000 136.200000 529.920000 136.300000 ;
      RECT 1.020000 135.320000 2.530000 136.200000 ;
      RECT 527.390000 135.120000 529.920000 136.200000 ;
      RECT 3.930000 135.120000 525.990000 136.200000 ;
      RECT 0.000000 135.120000 2.530000 135.320000 ;
      RECT 0.000000 133.480000 529.920000 135.120000 ;
      RECT 0.000000 133.250000 1.130000 133.480000 ;
      RECT 528.790000 132.400000 529.920000 133.480000 ;
      RECT 2.530000 132.400000 527.390000 133.480000 ;
      RECT 1.020000 132.400000 1.130000 133.250000 ;
      RECT 1.020000 132.270000 529.920000 132.400000 ;
      RECT 0.000000 130.760000 529.920000 132.270000 ;
      RECT 527.390000 129.680000 529.920000 130.760000 ;
      RECT 3.930000 129.680000 525.990000 130.760000 ;
      RECT 0.000000 129.680000 2.530000 130.760000 ;
      RECT 0.000000 129.590000 529.920000 129.680000 ;
      RECT 1.020000 128.610000 529.920000 129.590000 ;
      RECT 0.000000 128.040000 529.920000 128.610000 ;
      RECT 528.790000 126.960000 529.920000 128.040000 ;
      RECT 2.530000 126.960000 527.390000 128.040000 ;
      RECT 0.000000 126.960000 1.130000 128.040000 ;
      RECT 0.000000 126.540000 529.920000 126.960000 ;
      RECT 1.020000 125.560000 529.920000 126.540000 ;
      RECT 0.000000 125.320000 529.920000 125.560000 ;
      RECT 527.390000 124.240000 529.920000 125.320000 ;
      RECT 3.930000 124.240000 525.990000 125.320000 ;
      RECT 0.000000 124.240000 2.530000 125.320000 ;
      RECT 0.000000 122.880000 529.920000 124.240000 ;
      RECT 1.020000 122.600000 529.920000 122.880000 ;
      RECT 1.020000 121.900000 1.130000 122.600000 ;
      RECT 528.790000 121.520000 529.920000 122.600000 ;
      RECT 2.530000 121.520000 527.390000 122.600000 ;
      RECT 0.000000 121.520000 1.130000 121.900000 ;
      RECT 0.000000 119.880000 529.920000 121.520000 ;
      RECT 0.000000 119.830000 2.530000 119.880000 ;
      RECT 1.020000 118.850000 2.530000 119.830000 ;
      RECT 527.390000 118.800000 529.920000 119.880000 ;
      RECT 3.930000 118.800000 525.990000 119.880000 ;
      RECT 0.000000 118.800000 2.530000 118.850000 ;
      RECT 0.000000 117.160000 529.920000 118.800000 ;
      RECT 0.000000 116.170000 1.130000 117.160000 ;
      RECT 528.790000 116.080000 529.920000 117.160000 ;
      RECT 2.530000 116.080000 527.390000 117.160000 ;
      RECT 1.020000 116.080000 1.130000 116.170000 ;
      RECT 1.020000 115.190000 529.920000 116.080000 ;
      RECT 0.000000 114.440000 529.920000 115.190000 ;
      RECT 527.390000 113.360000 529.920000 114.440000 ;
      RECT 3.930000 113.360000 525.990000 114.440000 ;
      RECT 0.000000 113.360000 2.530000 114.440000 ;
      RECT 0.000000 113.120000 529.920000 113.360000 ;
      RECT 1.020000 112.140000 529.920000 113.120000 ;
      RECT 0.000000 111.720000 529.920000 112.140000 ;
      RECT 528.790000 110.640000 529.920000 111.720000 ;
      RECT 2.530000 110.640000 527.390000 111.720000 ;
      RECT 0.000000 110.640000 1.130000 111.720000 ;
      RECT 0.000000 109.460000 529.920000 110.640000 ;
      RECT 1.020000 109.000000 529.920000 109.460000 ;
      RECT 1.020000 108.480000 2.530000 109.000000 ;
      RECT 527.390000 107.920000 529.920000 109.000000 ;
      RECT 3.930000 107.920000 525.990000 109.000000 ;
      RECT 0.000000 107.920000 2.530000 108.480000 ;
      RECT 0.000000 106.410000 529.920000 107.920000 ;
      RECT 1.020000 106.280000 529.920000 106.410000 ;
      RECT 1.020000 105.430000 1.130000 106.280000 ;
      RECT 528.790000 105.200000 529.920000 106.280000 ;
      RECT 2.530000 105.200000 527.390000 106.280000 ;
      RECT 0.000000 105.200000 1.130000 105.430000 ;
      RECT 0.000000 103.560000 529.920000 105.200000 ;
      RECT 0.000000 102.750000 2.530000 103.560000 ;
      RECT 527.390000 102.480000 529.920000 103.560000 ;
      RECT 3.930000 102.480000 525.990000 103.560000 ;
      RECT 1.020000 102.480000 2.530000 102.750000 ;
      RECT 1.020000 101.770000 529.920000 102.480000 ;
      RECT 0.000000 100.840000 529.920000 101.770000 ;
      RECT 528.790000 99.760000 529.920000 100.840000 ;
      RECT 2.530000 99.760000 527.390000 100.840000 ;
      RECT 0.000000 99.760000 1.130000 100.840000 ;
      RECT 0.000000 99.700000 529.920000 99.760000 ;
      RECT 1.020000 98.720000 529.920000 99.700000 ;
      RECT 0.000000 98.120000 529.920000 98.720000 ;
      RECT 527.390000 97.040000 529.920000 98.120000 ;
      RECT 3.930000 97.040000 525.990000 98.120000 ;
      RECT 0.000000 97.040000 2.530000 98.120000 ;
      RECT 0.000000 96.040000 529.920000 97.040000 ;
      RECT 1.020000 95.400000 529.920000 96.040000 ;
      RECT 1.020000 95.060000 1.130000 95.400000 ;
      RECT 528.790000 94.320000 529.920000 95.400000 ;
      RECT 2.530000 94.320000 527.390000 95.400000 ;
      RECT 0.000000 94.320000 1.130000 95.060000 ;
      RECT 0.000000 92.990000 529.920000 94.320000 ;
      RECT 1.020000 92.680000 529.920000 92.990000 ;
      RECT 1.020000 92.010000 2.530000 92.680000 ;
      RECT 527.390000 91.600000 529.920000 92.680000 ;
      RECT 3.930000 91.600000 525.990000 92.680000 ;
      RECT 0.000000 91.600000 2.530000 92.010000 ;
      RECT 0.000000 89.960000 529.920000 91.600000 ;
      RECT 0.000000 89.330000 1.130000 89.960000 ;
      RECT 528.790000 88.880000 529.920000 89.960000 ;
      RECT 2.530000 88.880000 527.390000 89.960000 ;
      RECT 1.020000 88.880000 1.130000 89.330000 ;
      RECT 1.020000 88.350000 529.920000 88.880000 ;
      RECT 0.000000 87.240000 529.920000 88.350000 ;
      RECT 0.000000 86.280000 2.530000 87.240000 ;
      RECT 527.390000 86.160000 529.920000 87.240000 ;
      RECT 3.930000 86.160000 525.990000 87.240000 ;
      RECT 1.020000 86.160000 2.530000 86.280000 ;
      RECT 1.020000 85.300000 529.920000 86.160000 ;
      RECT 0.000000 84.520000 529.920000 85.300000 ;
      RECT 528.790000 83.440000 529.920000 84.520000 ;
      RECT 2.530000 83.440000 527.390000 84.520000 ;
      RECT 0.000000 83.440000 1.130000 84.520000 ;
      RECT 0.000000 82.620000 529.920000 83.440000 ;
      RECT 1.020000 81.800000 529.920000 82.620000 ;
      RECT 1.020000 81.640000 2.530000 81.800000 ;
      RECT 527.390000 80.720000 529.920000 81.800000 ;
      RECT 3.930000 80.720000 525.990000 81.800000 ;
      RECT 0.000000 80.720000 2.530000 81.640000 ;
      RECT 0.000000 79.570000 529.920000 80.720000 ;
      RECT 1.020000 79.080000 529.920000 79.570000 ;
      RECT 1.020000 78.590000 1.130000 79.080000 ;
      RECT 528.790000 78.000000 529.920000 79.080000 ;
      RECT 2.530000 78.000000 527.390000 79.080000 ;
      RECT 0.000000 78.000000 1.130000 78.590000 ;
      RECT 0.000000 76.360000 529.920000 78.000000 ;
      RECT 0.000000 75.910000 2.530000 76.360000 ;
      RECT 527.390000 75.280000 529.920000 76.360000 ;
      RECT 3.930000 75.280000 525.990000 76.360000 ;
      RECT 1.020000 75.280000 2.530000 75.910000 ;
      RECT 1.020000 74.930000 529.920000 75.280000 ;
      RECT 0.000000 73.640000 529.920000 74.930000 ;
      RECT 0.000000 72.860000 1.130000 73.640000 ;
      RECT 528.790000 72.560000 529.920000 73.640000 ;
      RECT 2.530000 72.560000 527.390000 73.640000 ;
      RECT 1.020000 72.560000 1.130000 72.860000 ;
      RECT 1.020000 71.880000 529.920000 72.560000 ;
      RECT 0.000000 70.920000 529.920000 71.880000 ;
      RECT 527.390000 69.840000 529.920000 70.920000 ;
      RECT 3.930000 69.840000 525.990000 70.920000 ;
      RECT 0.000000 69.840000 2.530000 70.920000 ;
      RECT 0.000000 69.200000 529.920000 69.840000 ;
      RECT 1.020000 68.220000 529.920000 69.200000 ;
      RECT 0.000000 68.200000 529.920000 68.220000 ;
      RECT 528.790000 67.120000 529.920000 68.200000 ;
      RECT 2.530000 67.120000 527.390000 68.200000 ;
      RECT 0.000000 67.120000 1.130000 68.200000 ;
      RECT 0.000000 66.150000 529.920000 67.120000 ;
      RECT 1.020000 65.480000 529.920000 66.150000 ;
      RECT 1.020000 65.170000 2.530000 65.480000 ;
      RECT 527.390000 64.400000 529.920000 65.480000 ;
      RECT 3.930000 64.400000 525.990000 65.480000 ;
      RECT 0.000000 64.400000 2.530000 65.170000 ;
      RECT 0.000000 62.760000 529.920000 64.400000 ;
      RECT 0.000000 62.490000 1.130000 62.760000 ;
      RECT 528.790000 61.680000 529.920000 62.760000 ;
      RECT 2.530000 61.680000 527.390000 62.760000 ;
      RECT 1.020000 61.680000 1.130000 62.490000 ;
      RECT 1.020000 61.510000 529.920000 61.680000 ;
      RECT 0.000000 60.040000 529.920000 61.510000 ;
      RECT 0.000000 59.440000 2.530000 60.040000 ;
      RECT 527.390000 58.960000 529.920000 60.040000 ;
      RECT 3.930000 58.960000 525.990000 60.040000 ;
      RECT 1.020000 58.960000 2.530000 59.440000 ;
      RECT 1.020000 58.460000 529.920000 58.960000 ;
      RECT 0.000000 57.320000 529.920000 58.460000 ;
      RECT 528.790000 56.240000 529.920000 57.320000 ;
      RECT 2.530000 56.240000 527.390000 57.320000 ;
      RECT 0.000000 56.240000 1.130000 57.320000 ;
      RECT 0.000000 55.780000 529.920000 56.240000 ;
      RECT 1.020000 54.800000 529.920000 55.780000 ;
      RECT 0.000000 54.600000 529.920000 54.800000 ;
      RECT 527.390000 53.520000 529.920000 54.600000 ;
      RECT 3.930000 53.520000 525.990000 54.600000 ;
      RECT 0.000000 53.520000 2.530000 54.600000 ;
      RECT 0.000000 52.730000 529.920000 53.520000 ;
      RECT 1.020000 51.880000 529.920000 52.730000 ;
      RECT 1.020000 51.750000 1.130000 51.880000 ;
      RECT 528.790000 50.800000 529.920000 51.880000 ;
      RECT 2.530000 50.800000 527.390000 51.880000 ;
      RECT 0.000000 50.800000 1.130000 51.750000 ;
      RECT 0.000000 49.160000 529.920000 50.800000 ;
      RECT 0.000000 49.070000 2.530000 49.160000 ;
      RECT 1.020000 48.090000 2.530000 49.070000 ;
      RECT 527.390000 48.080000 529.920000 49.160000 ;
      RECT 3.930000 48.080000 525.990000 49.160000 ;
      RECT 0.000000 48.080000 2.530000 48.090000 ;
      RECT 0.000000 46.440000 529.920000 48.080000 ;
      RECT 0.000000 46.020000 1.130000 46.440000 ;
      RECT 528.790000 45.360000 529.920000 46.440000 ;
      RECT 2.530000 45.360000 527.390000 46.440000 ;
      RECT 1.020000 45.360000 1.130000 46.020000 ;
      RECT 1.020000 45.040000 529.920000 45.360000 ;
      RECT 0.000000 43.720000 529.920000 45.040000 ;
      RECT 527.390000 42.640000 529.920000 43.720000 ;
      RECT 3.930000 42.640000 525.990000 43.720000 ;
      RECT 0.000000 42.640000 2.530000 43.720000 ;
      RECT 0.000000 42.360000 529.920000 42.640000 ;
      RECT 1.020000 41.380000 529.920000 42.360000 ;
      RECT 0.000000 41.000000 529.920000 41.380000 ;
      RECT 528.790000 39.920000 529.920000 41.000000 ;
      RECT 2.530000 39.920000 527.390000 41.000000 ;
      RECT 0.000000 39.920000 1.130000 41.000000 ;
      RECT 0.000000 39.310000 529.920000 39.920000 ;
      RECT 1.020000 38.330000 529.920000 39.310000 ;
      RECT 0.000000 38.280000 529.920000 38.330000 ;
      RECT 527.390000 37.200000 529.920000 38.280000 ;
      RECT 3.930000 37.200000 525.990000 38.280000 ;
      RECT 0.000000 37.200000 2.530000 38.280000 ;
      RECT 0.000000 35.650000 529.920000 37.200000 ;
      RECT 1.020000 35.560000 529.920000 35.650000 ;
      RECT 1.020000 34.670000 1.130000 35.560000 ;
      RECT 528.790000 34.480000 529.920000 35.560000 ;
      RECT 2.530000 34.480000 527.390000 35.560000 ;
      RECT 0.000000 34.480000 1.130000 34.670000 ;
      RECT 0.000000 32.840000 529.920000 34.480000 ;
      RECT 0.000000 32.600000 2.530000 32.840000 ;
      RECT 527.390000 31.760000 529.920000 32.840000 ;
      RECT 3.930000 31.760000 525.990000 32.840000 ;
      RECT 1.020000 31.760000 2.530000 32.600000 ;
      RECT 1.020000 31.620000 529.920000 31.760000 ;
      RECT 0.000000 30.120000 529.920000 31.620000 ;
      RECT 528.790000 29.040000 529.920000 30.120000 ;
      RECT 2.530000 29.040000 527.390000 30.120000 ;
      RECT 0.000000 29.040000 1.130000 30.120000 ;
      RECT 0.000000 28.940000 529.920000 29.040000 ;
      RECT 1.020000 27.960000 529.920000 28.940000 ;
      RECT 0.000000 27.400000 529.920000 27.960000 ;
      RECT 527.390000 26.320000 529.920000 27.400000 ;
      RECT 3.930000 26.320000 525.990000 27.400000 ;
      RECT 0.000000 26.320000 2.530000 27.400000 ;
      RECT 0.000000 25.890000 529.920000 26.320000 ;
      RECT 1.020000 24.910000 529.920000 25.890000 ;
      RECT 0.000000 24.680000 529.920000 24.910000 ;
      RECT 528.790000 23.600000 529.920000 24.680000 ;
      RECT 2.530000 23.600000 527.390000 24.680000 ;
      RECT 0.000000 23.600000 1.130000 24.680000 ;
      RECT 0.000000 22.230000 529.920000 23.600000 ;
      RECT 1.020000 21.960000 529.920000 22.230000 ;
      RECT 1.020000 21.250000 2.530000 21.960000 ;
      RECT 527.390000 20.880000 529.920000 21.960000 ;
      RECT 3.930000 20.880000 525.990000 21.960000 ;
      RECT 0.000000 20.880000 2.530000 21.250000 ;
      RECT 0.000000 19.240000 529.920000 20.880000 ;
      RECT 0.000000 19.180000 1.130000 19.240000 ;
      RECT 1.020000 18.200000 1.130000 19.180000 ;
      RECT 528.790000 18.160000 529.920000 19.240000 ;
      RECT 2.530000 18.160000 527.390000 19.240000 ;
      RECT 0.000000 18.160000 1.130000 18.200000 ;
      RECT 0.000000 16.520000 529.920000 18.160000 ;
      RECT 0.000000 15.520000 2.530000 16.520000 ;
      RECT 527.390000 15.440000 529.920000 16.520000 ;
      RECT 3.930000 15.440000 525.990000 16.520000 ;
      RECT 1.020000 15.440000 2.530000 15.520000 ;
      RECT 1.020000 14.540000 529.920000 15.440000 ;
      RECT 0.000000 13.800000 529.920000 14.540000 ;
      RECT 528.790000 12.720000 529.920000 13.800000 ;
      RECT 2.530000 12.720000 527.390000 13.800000 ;
      RECT 0.000000 12.720000 1.130000 13.800000 ;
      RECT 0.000000 12.470000 529.920000 12.720000 ;
      RECT 1.020000 11.490000 529.920000 12.470000 ;
      RECT 0.000000 11.080000 529.920000 11.490000 ;
      RECT 527.390000 10.000000 529.920000 11.080000 ;
      RECT 3.930000 10.000000 525.990000 11.080000 ;
      RECT 0.000000 10.000000 2.530000 11.080000 ;
      RECT 0.000000 8.810000 529.920000 10.000000 ;
      RECT 1.020000 8.360000 529.920000 8.810000 ;
      RECT 1.020000 7.830000 1.130000 8.360000 ;
      RECT 528.790000 7.280000 529.920000 8.360000 ;
      RECT 2.530000 7.280000 527.390000 8.360000 ;
      RECT 0.000000 7.280000 1.130000 7.830000 ;
      RECT 0.000000 5.760000 529.920000 7.280000 ;
      RECT 1.020000 5.640000 529.920000 5.760000 ;
      RECT 1.020000 4.780000 2.530000 5.640000 ;
      RECT 527.390000 4.560000 529.920000 5.640000 ;
      RECT 3.930000 4.560000 525.990000 5.640000 ;
      RECT 0.000000 4.560000 2.530000 4.780000 ;
      RECT 0.000000 3.950000 529.920000 4.560000 ;
      RECT 0.000000 2.550000 2.530000 3.950000 ;
      RECT 0.000000 1.150000 1.130000 2.550000 ;
      RECT 0.000000 0.000000 529.920000 1.150000 ;
    LAYER met4 ;
      RECT 528.790000 0.000000 529.920000 420.240000 ;
      RECT 3.930000 0.000000 525.990000 420.240000 ;
      RECT 0.000000 0.000000 1.130000 420.240000 ;
  END
END BlockRAM_1KB

END LIBRARY
