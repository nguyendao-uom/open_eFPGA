##
## LEF for PtnCells ;
## created by Innovus v19.11-s128_1 on Fri Dec  3 16:33:23 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO ibex_core
  CLASS BLOCK ;
  SIZE 550.160000 BY 549.780000 ;
  FOREIGN ibex_core 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.4511 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5585 LAYER met3  ;
    ANTENNAMAXAREACAR 59.5278 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 300.108 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 9.840000 550.160000 10.220000 ;
    END
  END clk_i
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8765 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.328 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 13.2483 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 67.5273 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 137.626 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 737.752 LAYER met4  ;
    ANTENNAGATEAREA 3.327 LAYER met4  ;
    ANTENNAMAXAREACAR 125.647 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 666.741 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.854141 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 11.670000 550.160000 12.050000 ;
    END
  END rst_ni
  PIN test_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 22.8556 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 108.476 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 14.110000 550.160000 14.490000 ;
    END
  END test_en_i
  PIN core_id_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.894 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.704 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 53.159 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 278.982 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 16.550000 550.160000 16.930000 ;
    END
  END core_id_i[3]
  PIN core_id_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.5112 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 43.7699 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 235.261 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 18.990000 550.160000 19.370000 ;
    END
  END core_id_i[2]
  PIN core_id_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.351 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 99.9897 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 507.41 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 20.820000 550.160000 21.200000 ;
    END
  END core_id_i[1]
  PIN core_id_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 21.1683 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 102.044 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 23.260000 550.160000 23.640000 ;
    END
  END core_id_i[0]
  PIN cluster_id_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.815 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 128.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 23.8261 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 124.594 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 25.700000 550.160000 26.080000 ;
    END
  END cluster_id_i[5]
  PIN cluster_id_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.2786 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 45.1752 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 246.299 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 28.140000 550.160000 28.520000 ;
    END
  END cluster_id_i[4]
  PIN cluster_id_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.0428 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 156.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 60.4949 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 314.683 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 29.970000 550.160000 30.350000 ;
    END
  END cluster_id_i[3]
  PIN cluster_id_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.224 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 27.0802 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 134.913 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 32.410000 550.160000 32.790000 ;
    END
  END cluster_id_i[2]
  PIN cluster_id_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 73.9531 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 396.489 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 34.850000 550.160000 35.230000 ;
    END
  END cluster_id_i[1]
  PIN cluster_id_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.1398 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 37.66 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 192.113 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 37.290000 550.160000 37.670000 ;
    END
  END cluster_id_i[0]
  PIN boot_addr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.9006 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 52.6554 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 282.24 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 87.5436 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 462.085 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.423165 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 39.120000 550.160000 39.500000 ;
    END
  END boot_addr_i[31]
  PIN boot_addr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.1356 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 166.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 46.2348 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 247.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 74.2632 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 391.897 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.315421 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 41.560000 550.160000 41.940000 ;
    END
  END boot_addr_i[30]
  PIN boot_addr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 38.8666 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 207.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.1938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 241.504 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 96.904 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 495.347 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.536761 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 44.000000 550.160000 44.380000 ;
    END
  END boot_addr_i[29]
  PIN boot_addr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.6566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 174.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.1368 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 241.2 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 94.7908 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 499.228 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.536761 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 46.440000 550.160000 46.820000 ;
    END
  END boot_addr_i[28]
  PIN boot_addr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.2126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 39.0186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 209.04 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 74.4092 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 386.319 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.536761 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 48.270000 550.160000 48.650000 ;
    END
  END boot_addr_i[27]
  PIN boot_addr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.5294 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.9006 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 245.744 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 83.405 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 434.584 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.536761 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 50.710000 550.160000 51.090000 ;
    END
  END boot_addr_i[26]
  PIN boot_addr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.1456 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 128.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 44.5806 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 238.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 89.5696 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 465.911 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.536761 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 53.150000 550.160000 53.530000 ;
    END
  END boot_addr_i[25]
  PIN boot_addr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.9854 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.5086 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 222.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 88.7652 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 459.027 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.536761 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 55.590000 550.160000 55.970000 ;
    END
  END boot_addr_i[24]
  PIN boot_addr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4586 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.9292 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 225.504 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 81.5188 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 426.237 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.536761 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 57.420000 550.160000 57.800000 ;
    END
  END boot_addr_i[23]
  PIN boot_addr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 42.7744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 230.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 26.0718 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 118.232 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.536761 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 59.860000 550.160000 60.240000 ;
    END
  END boot_addr_i[22]
  PIN boot_addr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.152 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 30.3294 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 163.168 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 83.1414 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 434.359 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.536761 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 62.300000 550.160000 62.680000 ;
    END
  END boot_addr_i[21]
  PIN boot_addr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 38.1016 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 203.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 37.3476 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 200.128 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 84.7372 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 432.45 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.536761 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 64.740000 550.160000 65.120000 ;
    END
  END boot_addr_i[20]
  PIN boot_addr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 43.1896 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 230.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 39.6078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 211.712 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 77.9352 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 397.488 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.536761 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 66.570000 550.160000 66.950000 ;
    END
  END boot_addr_i[19]
  PIN boot_addr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.554 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 169.224 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met3  ;
    ANTENNAMAXAREACAR 72.3799 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 370.251 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.472349 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 69.010000 550.160000 69.390000 ;
    END
  END boot_addr_i[18]
  PIN boot_addr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.4586 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 189.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.3748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 173.136 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 72.8012 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 374.325 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.536761 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 71.450000 550.160000 71.830000 ;
    END
  END boot_addr_i[17]
  PIN boot_addr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 34.0816 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 181.76 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.2187 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 241.632 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 97.6211 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 509.784 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 73.890000 550.160000 74.270000 ;
    END
  END boot_addr_i[16]
  PIN boot_addr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 28.7956 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 153.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 36.0348 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 192.656 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 78.1268 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 402.934 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.536761 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 75.720000 550.160000 76.100000 ;
    END
  END boot_addr_i[15]
  PIN boot_addr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 30.8416 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 164.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 28.8738 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 154.464 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 72.6183 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 366.714 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.536761 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 78.160000 550.160000 78.540000 ;
    END
  END boot_addr_i[14]
  PIN boot_addr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.8956 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 148.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 36.6168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 195.76 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 66.8234 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 345.989 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.536761 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 80.600000 550.160000 80.980000 ;
    END
  END boot_addr_i[13]
  PIN boot_addr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.5246 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125.456 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 34.5078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 184.512 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 56.9486 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 298.133 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.315421 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 83.040000 550.160000 83.420000 ;
    END
  END boot_addr_i[12]
  PIN boot_addr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1756 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 37.4508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 200.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 80.4642 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 426.642 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.315421 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 84.870000 550.160000 85.250000 ;
    END
  END boot_addr_i[11]
  PIN boot_addr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7774 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 32.5094 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 169.497 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.315421 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 87.310000 550.160000 87.690000 ;
    END
  END boot_addr_i[10]
  PIN boot_addr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6246 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.5656 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 174.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 66.6684 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 348.945 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.423165 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 89.750000 550.160000 90.130000 ;
    END
  END boot_addr_i[9]
  PIN boot_addr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.6146 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 38.9706 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 208.784 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 71.6259 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 382.522 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 92.190000 550.160000 92.570000 ;
    END
  END boot_addr_i[8]
  PIN boot_addr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.1292 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.488 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 57.5051 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 303.2 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 94.630000 550.160000 95.010000 ;
    END
  END boot_addr_i[7]
  PIN boot_addr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.1374 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 52.2006 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 272.384 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 96.460000 550.160000 96.840000 ;
    END
  END boot_addr_i[6]
  PIN boot_addr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.8626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.4336 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 18.545 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 98.804 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 98.900000 550.160000 99.280000 ;
    END
  END boot_addr_i[5]
  PIN boot_addr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.7972 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 135.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 13.2145 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 70.5414 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 101.340000 550.160000 101.720000 ;
    END
  END boot_addr_i[4]
  PIN boot_addr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 39.2352 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 192.057 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 103.780000 550.160000 104.160000 ;
    END
  END boot_addr_i[3]
  PIN boot_addr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.1948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.112 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 87.0085 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 455.547 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 105.610000 550.160000 105.990000 ;
    END
  END boot_addr_i[2]
  PIN boot_addr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.8888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 63.9188 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 328.23 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 108.050000 550.160000 108.430000 ;
    END
  END boot_addr_i[1]
  PIN boot_addr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.07 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 21.063 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 109.859 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 110.490000 550.160000 110.870000 ;
    END
  END boot_addr_i[0]
  PIN instr_req_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 112.930000 550.160000 113.310000 ;
    END
  END instr_req_o
  PIN instr_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.888 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met3  ;
    ANTENNAMAXAREACAR 13.9801 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 54.246 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.335662 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 114.760000 550.160000 115.140000 ;
    END
  END instr_gnt_i
  PIN instr_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met3  ;
    ANTENNAMAXAREACAR 7.6172 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 36.5193 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.453993 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 117.200000 550.160000 117.580000 ;
    END
  END instr_rvalid_i
  PIN instr_addr_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 33.5694 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 179.032 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 119.640000 550.160000 120.020000 ;
    END
  END instr_addr_o[31]
  PIN instr_addr_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 35.2134 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 187.8 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 122.080000 550.160000 122.460000 ;
    END
  END instr_addr_o[30]
  PIN instr_addr_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 38.3004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 204.264 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 123.910000 550.160000 124.290000 ;
    END
  END instr_addr_o[29]
  PIN instr_addr_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 163.816 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 126.350000 550.160000 126.730000 ;
    END
  END instr_addr_o[28]
  PIN instr_addr_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 31.4382 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 168.136 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 128.790000 550.160000 129.170000 ;
    END
  END instr_addr_o[27]
  PIN instr_addr_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.7176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 131.230000 550.160000 131.610000 ;
    END
  END instr_addr_o[26]
  PIN instr_addr_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 40.0846 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 213.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.9378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.472 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 133.060000 550.160000 133.440000 ;
    END
  END instr_addr_o[25]
  PIN instr_addr_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 39.8274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 212.408 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 135.500000 550.160000 135.880000 ;
    END
  END instr_addr_o[24]
  PIN instr_addr_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 42.9954 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 229.304 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 137.940000 550.160000 138.320000 ;
    END
  END instr_addr_o[23]
  PIN instr_addr_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.7026 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 140.380000 550.160000 140.760000 ;
    END
  END instr_addr_o[22]
  PIN instr_addr_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 36.9714 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 197.176 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 142.210000 550.160000 142.590000 ;
    END
  END instr_addr_o[21]
  PIN instr_addr_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.5346 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.6166 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.896 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 144.650000 550.160000 145.030000 ;
    END
  END instr_addr_o[20]
  PIN instr_addr_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.6152 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.08 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 147.090000 550.160000 147.470000 ;
    END
  END instr_addr_o[19]
  PIN instr_addr_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.9262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 144.072 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 149.530000 550.160000 149.910000 ;
    END
  END instr_addr_o[18]
  PIN instr_addr_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.482 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.84 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 151.360000 550.160000 151.740000 ;
    END
  END instr_addr_o[17]
  PIN instr_addr_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.4426 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 153.800000 550.160000 154.180000 ;
    END
  END instr_addr_o[16]
  PIN instr_addr_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 156.240000 550.160000 156.620000 ;
    END
  END instr_addr_o[15]
  PIN instr_addr_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 158.680000 550.160000 159.060000 ;
    END
  END instr_addr_o[14]
  PIN instr_addr_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.4124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.528 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 160.510000 550.160000 160.890000 ;
    END
  END instr_addr_o[13]
  PIN instr_addr_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.4144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 162.950000 550.160000 163.330000 ;
    END
  END instr_addr_o[12]
  PIN instr_addr_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 165.390000 550.160000 165.770000 ;
    END
  END instr_addr_o[11]
  PIN instr_addr_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.9414 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.016 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 167.830000 550.160000 168.210000 ;
    END
  END instr_addr_o[10]
  PIN instr_addr_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 170.270000 550.160000 170.650000 ;
    END
  END instr_addr_o[9]
  PIN instr_addr_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.3524 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.208 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 172.100000 550.160000 172.480000 ;
    END
  END instr_addr_o[8]
  PIN instr_addr_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.4124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.528 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 174.540000 550.160000 174.920000 ;
    END
  END instr_addr_o[7]
  PIN instr_addr_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 176.980000 550.160000 177.360000 ;
    END
  END instr_addr_o[6]
  PIN instr_addr_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 179.420000 550.160000 179.800000 ;
    END
  END instr_addr_o[5]
  PIN instr_addr_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 181.250000 550.160000 181.630000 ;
    END
  END instr_addr_o[4]
  PIN instr_addr_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 183.690000 550.160000 184.070000 ;
    END
  END instr_addr_o[3]
  PIN instr_addr_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 186.130000 550.160000 186.510000 ;
    END
  END instr_addr_o[2]
  PIN instr_addr_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 188.570000 550.160000 188.950000 ;
    END
  END instr_addr_o[1]
  PIN instr_addr_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.8034 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 190.400000 550.160000 190.780000 ;
    END
  END instr_addr_o[0]
  PIN instr_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9524 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.7788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 53.3102 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 266.651 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.14868 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 192.840000 550.160000 193.220000 ;
    END
  END instr_rdata_i[31]
  PIN instr_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.5686 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.024 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.1878 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 113.472 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 98.3118 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 500.085 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.798148 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 195.280000 550.160000 195.660000 ;
    END
  END instr_rdata_i[30]
  PIN instr_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met3  ;
    ANTENNAMAXAREACAR 30.8484 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 141.957 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.513757 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 197.720000 550.160000 198.100000 ;
    END
  END instr_rdata_i[29]
  PIN instr_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.4983 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.064 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met3  ;
    ANTENNAMAXAREACAR 103.731 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 520.511 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 199.550000 550.160000 199.930000 ;
    END
  END instr_rdata_i[28]
  PIN instr_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.824 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met3  ;
    ANTENNAMAXAREACAR 62.2437 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 308.256 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 201.990000 550.160000 202.370000 ;
    END
  END instr_rdata_i[27]
  PIN instr_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met3  ;
    ANTENNAMAXAREACAR 38.0386 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 178.366 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.513757 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 204.430000 550.160000 204.810000 ;
    END
  END instr_rdata_i[26]
  PIN instr_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.096 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met3  ;
    ANTENNAMAXAREACAR 98.3694 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.31 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 206.870000 550.160000 207.250000 ;
    END
  END instr_rdata_i[25]
  PIN instr_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.7458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 68.448 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 76.0602 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 385.567 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32725 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 208.700000 550.160000 209.080000 ;
    END
  END instr_rdata_i[24]
  PIN instr_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met3  ;
    ANTENNAMAXAREACAR 74.1036 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 356.406 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.692328 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 211.140000 550.160000 211.520000 ;
    END
  END instr_rdata_i[23]
  PIN instr_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.2911 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.68 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met3  ;
    ANTENNAMAXAREACAR 74.6472 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 372.171 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 213.580000 550.160000 213.960000 ;
    END
  END instr_rdata_i[22]
  PIN instr_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4096 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met3  ;
    ANTENNAMAXAREACAR 143.854 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 720.422 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 216.020000 550.160000 216.400000 ;
    END
  END instr_rdata_i[21]
  PIN instr_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met3  ;
    ANTENNAMAXAREACAR 32.6571 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 151.065 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.513757 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 217.850000 550.160000 218.230000 ;
    END
  END instr_rdata_i[20]
  PIN instr_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met3  ;
    ANTENNAMAXAREACAR 66.3041 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 317.647 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.692328 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 220.290000 550.160000 220.670000 ;
    END
  END instr_rdata_i[19]
  PIN instr_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met3  ;
    ANTENNAMAXAREACAR 61.9165 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 293.897 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.870899 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 222.730000 550.160000 223.110000 ;
    END
  END instr_rdata_i[18]
  PIN instr_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.4544 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.3558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.368 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 79.7427 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 406.224 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.851058 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 225.170000 550.160000 225.550000 ;
    END
  END instr_rdata_i[17]
  PIN instr_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.3382 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.936 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met3  ;
    ANTENNAMAXAREACAR 59.6134 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 297.251 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.513757 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 227.000000 550.160000 227.380000 ;
    END
  END instr_rdata_i[16]
  PIN instr_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.2556 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.04 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9774 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 57.5488 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 293.595 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 229.440000 550.160000 229.820000 ;
    END
  END instr_rdata_i[15]
  PIN instr_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.42 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 132.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met3  ;
    ANTENNAMAXAREACAR 77.9623 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 402.475 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 231.880000 550.160000 232.260000 ;
    END
  END instr_rdata_i[14]
  PIN instr_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0472 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.384 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met3  ;
    ANTENNAMAXAREACAR 58.0948 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 279.254 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.513757 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 234.320000 550.160000 234.700000 ;
    END
  END instr_rdata_i[13]
  PIN instr_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.3258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 48.2302 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 237.05 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.619577 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 236.150000 550.160000 236.530000 ;
    END
  END instr_rdata_i[12]
  PIN instr_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.044 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met3  ;
    ANTENNAMAXAREACAR 87.4475 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 443.284 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.692328 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 238.590000 550.160000 238.970000 ;
    END
  END instr_rdata_i[11]
  PIN instr_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.8296 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 128.032 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met3  ;
    ANTENNAMAXAREACAR 83.044 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 421.745 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 241.030000 550.160000 241.410000 ;
    END
  END instr_rdata_i[10]
  PIN instr_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.3562 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 95.384 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met3  ;
    ANTENNAMAXAREACAR 88.6631 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 453.717 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.394709 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 243.470000 550.160000 243.850000 ;
    END
  END instr_rdata_i[9]
  PIN instr_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.6064 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.664 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 62.0623 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 329.44 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.67778 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 245.910000 550.160000 246.290000 ;
    END
  END instr_rdata_i[8]
  PIN instr_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.9475 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 45.9425 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 232.603 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 247.740000 550.160000 248.120000 ;
    END
  END instr_rdata_i[7]
  PIN instr_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.0832 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.0204 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 113.52 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 114.921 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 601.489 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.831217 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 250.180000 550.160000 250.560000 ;
    END
  END instr_rdata_i[6]
  PIN instr_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met3  ;
    ANTENNAMAXAREACAR 33.0097 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 151.415 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.513757 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 252.620000 550.160000 253.000000 ;
    END
  END instr_rdata_i[5]
  PIN instr_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.3534 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.816 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 88.4306 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 440.126 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.97672 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 255.060000 550.160000 255.440000 ;
    END
  END instr_rdata_i[4]
  PIN instr_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.4738 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 148.4 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 78.0968 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 405.891 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 256.890000 550.160000 257.270000 ;
    END
  END instr_rdata_i[3]
  PIN instr_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.1172 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 94.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2954 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 58.8094 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 302.302 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.831217 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 259.330000 550.160000 259.710000 ;
    END
  END instr_rdata_i[2]
  PIN instr_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.3014 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 121.288 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met3  ;
    ANTENNAMAXAREACAR 91.1393 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 466.042 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 261.770000 550.160000 262.150000 ;
    END
  END instr_rdata_i[1]
  PIN instr_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.1354 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 25.6518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 137.28 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met4  ;
    ANTENNAMAXAREACAR 121.764 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 622.985 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.798148 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 264.210000 550.160000 264.590000 ;
    END
  END instr_rdata_i[0]
  PIN data_req_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 266.040000 550.160000 266.420000 ;
    END
  END data_req_o
  PIN data_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9796 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.3778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 93.152 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0555 LAYER met4  ;
    ANTENNAMAXAREACAR 24.7643 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 117.681 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.618965 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 268.480000 550.160000 268.860000 ;
    END
  END data_gnt_i
  PIN data_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7136 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.0244 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 140.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 8.811 LAYER met4  ;
    ANTENNAMAXAREACAR 36.9437 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 183.562 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 270.920000 550.160000 271.300000 ;
    END
  END data_rvalid_i
  PIN data_we_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.5594 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.312 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 273.360000 550.160000 273.740000 ;
    END
  END data_we_o
  PIN data_be_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.4804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.224 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 275.190000 550.160000 275.570000 ;
    END
  END data_be_o[3]
  PIN data_be_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.4124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.528 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 277.630000 550.160000 278.010000 ;
    END
  END data_be_o[2]
  PIN data_be_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 280.070000 550.160000 280.450000 ;
    END
  END data_be_o[1]
  PIN data_be_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.6524 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.808 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 282.510000 550.160000 282.890000 ;
    END
  END data_be_o[0]
  PIN data_addr_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.3924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 162.088 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 284.340000 550.160000 284.720000 ;
    END
  END data_addr_o[31]
  PIN data_addr_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 27.8634 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 148.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 286.780000 550.160000 287.160000 ;
    END
  END data_addr_o[30]
  PIN data_addr_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.9762 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 165.672 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 289.220000 550.160000 289.600000 ;
    END
  END data_addr_o[29]
  PIN data_addr_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.2476 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.6218 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 41.12 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 291.660000 550.160000 292.040000 ;
    END
  END data_addr_o[28]
  PIN data_addr_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0036 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.7822 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.72 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 293.490000 550.160000 293.870000 ;
    END
  END data_addr_o[27]
  PIN data_addr_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 33.1842 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 177.448 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 295.930000 550.160000 296.310000 ;
    END
  END data_addr_o[26]
  PIN data_addr_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.6296 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.632 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 298.370000 550.160000 298.750000 ;
    END
  END data_addr_o[25]
  PIN data_addr_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 47.9154 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 255.544 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 300.810000 550.160000 301.190000 ;
    END
  END data_addr_o[24]
  PIN data_addr_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.7326 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.888 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 302.640000 550.160000 303.020000 ;
    END
  END data_addr_o[23]
  PIN data_addr_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 23.1582 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.976 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 305.080000 550.160000 305.460000 ;
    END
  END data_addr_o[22]
  PIN data_addr_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2456 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.8256 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.344 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 307.520000 550.160000 307.900000 ;
    END
  END data_addr_o[21]
  PIN data_addr_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 40.6576 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 216.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.4966 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.256 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 309.960000 550.160000 310.340000 ;
    END
  END data_addr_o[20]
  PIN data_addr_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5326 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.2082 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 226.992 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 311.790000 550.160000 312.170000 ;
    END
  END data_addr_o[19]
  PIN data_addr_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 38.3994 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 204.792 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 314.230000 550.160000 314.610000 ;
    END
  END data_addr_o[18]
  PIN data_addr_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2776 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 316.670000 550.160000 317.050000 ;
    END
  END data_addr_o[17]
  PIN data_addr_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.3924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 103.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.2908 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.688 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 319.110000 550.160000 319.490000 ;
    END
  END data_addr_o[16]
  PIN data_addr_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 321.550000 550.160000 321.930000 ;
    END
  END data_addr_o[15]
  PIN data_addr_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.2152 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 323.380000 550.160000 323.760000 ;
    END
  END data_addr_o[14]
  PIN data_addr_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0746 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.056 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.3538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 45.024 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 325.820000 550.160000 326.200000 ;
    END
  END data_addr_o[13]
  PIN data_addr_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.496 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.1086 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 81.52 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 328.260000 550.160000 328.640000 ;
    END
  END data_addr_o[12]
  PIN data_addr_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.2176 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 60.768 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 330.700000 550.160000 331.080000 ;
    END
  END data_addr_o[11]
  PIN data_addr_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.3016 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.4888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 77.744 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 332.530000 550.160000 332.910000 ;
    END
  END data_addr_o[10]
  PIN data_addr_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.5844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.112 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 334.970000 550.160000 335.350000 ;
    END
  END data_addr_o[9]
  PIN data_addr_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.8604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.584 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 337.410000 550.160000 337.790000 ;
    END
  END data_addr_o[8]
  PIN data_addr_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 339.850000 550.160000 340.230000 ;
    END
  END data_addr_o[7]
  PIN data_addr_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.496 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.4238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.064 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 341.680000 550.160000 342.060000 ;
    END
  END data_addr_o[6]
  PIN data_addr_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.6634 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.2 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 344.120000 550.160000 344.500000 ;
    END
  END data_addr_o[5]
  PIN data_addr_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 346.560000 550.160000 346.940000 ;
    END
  END data_addr_o[4]
  PIN data_addr_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 349.000000 550.160000 349.380000 ;
    END
  END data_addr_o[3]
  PIN data_addr_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.4464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.376 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 350.830000 550.160000 351.210000 ;
    END
  END data_addr_o[2]
  PIN data_addr_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.8944 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.432 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 353.270000 550.160000 353.650000 ;
    END
  END data_addr_o[1]
  PIN data_addr_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 355.710000 550.160000 356.090000 ;
    END
  END data_addr_o[0]
  PIN data_wdata_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 358.150000 550.160000 358.530000 ;
    END
  END data_wdata_o[31]
  PIN data_wdata_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 359.980000 550.160000 360.360000 ;
    END
  END data_wdata_o[30]
  PIN data_wdata_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.4234 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 362.420000 550.160000 362.800000 ;
    END
  END data_wdata_o[29]
  PIN data_wdata_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.2554 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.024 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 364.860000 550.160000 365.240000 ;
    END
  END data_wdata_o[28]
  PIN data_wdata_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.2514 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.336 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 367.300000 550.160000 367.680000 ;
    END
  END data_wdata_o[27]
  PIN data_wdata_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 369.130000 550.160000 369.510000 ;
    END
  END data_wdata_o[26]
  PIN data_wdata_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 371.570000 550.160000 371.950000 ;
    END
  END data_wdata_o[25]
  PIN data_wdata_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 374.010000 550.160000 374.390000 ;
    END
  END data_wdata_o[24]
  PIN data_wdata_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 376.450000 550.160000 376.830000 ;
    END
  END data_wdata_o[23]
  PIN data_wdata_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 378.280000 550.160000 378.660000 ;
    END
  END data_wdata_o[22]
  PIN data_wdata_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.0664 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.016 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 380.720000 550.160000 381.100000 ;
    END
  END data_wdata_o[21]
  PIN data_wdata_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.8164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.016 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 383.160000 550.160000 383.540000 ;
    END
  END data_wdata_o[20]
  PIN data_wdata_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 385.600000 550.160000 385.980000 ;
    END
  END data_wdata_o[19]
  PIN data_wdata_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 387.430000 550.160000 387.810000 ;
    END
  END data_wdata_o[18]
  PIN data_wdata_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 389.870000 550.160000 390.250000 ;
    END
  END data_wdata_o[17]
  PIN data_wdata_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 392.310000 550.160000 392.690000 ;
    END
  END data_wdata_o[16]
  PIN data_wdata_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.7944 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.232 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 394.750000 550.160000 395.130000 ;
    END
  END data_wdata_o[15]
  PIN data_wdata_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.1384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.4 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 397.190000 550.160000 397.570000 ;
    END
  END data_wdata_o[14]
  PIN data_wdata_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 399.020000 550.160000 399.400000 ;
    END
  END data_wdata_o[13]
  PIN data_wdata_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 401.460000 550.160000 401.840000 ;
    END
  END data_wdata_o[12]
  PIN data_wdata_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 403.900000 550.160000 404.280000 ;
    END
  END data_wdata_o[11]
  PIN data_wdata_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 406.340000 550.160000 406.720000 ;
    END
  END data_wdata_o[10]
  PIN data_wdata_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.4524 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.408 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 408.170000 550.160000 408.550000 ;
    END
  END data_wdata_o[9]
  PIN data_wdata_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.2964 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.576 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 410.610000 550.160000 410.990000 ;
    END
  END data_wdata_o[8]
  PIN data_wdata_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.7004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.064 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 413.050000 550.160000 413.430000 ;
    END
  END data_wdata_o[7]
  PIN data_wdata_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 415.490000 550.160000 415.870000 ;
    END
  END data_wdata_o[6]
  PIN data_wdata_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 417.320000 550.160000 417.700000 ;
    END
  END data_wdata_o[5]
  PIN data_wdata_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 419.760000 550.160000 420.140000 ;
    END
  END data_wdata_o[4]
  PIN data_wdata_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.0034 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 106.68 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 422.200000 550.160000 422.580000 ;
    END
  END data_wdata_o[3]
  PIN data_wdata_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.8284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 111.08 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 424.640000 550.160000 425.020000 ;
    END
  END data_wdata_o[2]
  PIN data_wdata_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 426.470000 550.160000 426.850000 ;
    END
  END data_wdata_o[1]
  PIN data_wdata_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 428.910000 550.160000 429.290000 ;
    END
  END data_wdata_o[0]
  PIN data_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9906 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.7308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 52.368 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 32.7015 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 152.988 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.515032 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 431.350000 550.160000 431.730000 ;
    END
  END data_rdata_i[31]
  PIN data_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.5153 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.872 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 24.0725 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 127.958 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.7068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 36.24 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 33.0508 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 176.472 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 433.790000 550.160000 434.170000 ;
    END
  END data_rdata_i[30]
  PIN data_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6864 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.656 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 18.2098 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 88.5936 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.640055 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 435.620000 550.160000 436.000000 ;
    END
  END data_rdata_i[29]
  PIN data_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.8988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 36.9819 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 174.752 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 438.060000 550.160000 438.440000 ;
    END
  END data_rdata_i[28]
  PIN data_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.16535 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.608 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 18.9185 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 98.7849 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.346263 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.2436 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.24 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 105.637 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 547.367 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.67778 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 440.500000 550.160000 440.880000 ;
    END
  END data_rdata_i[27]
  PIN data_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.5912 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.952 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 29.0936 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 133.739 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.477381 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 442.940000 550.160000 443.320000 ;
    END
  END data_rdata_i[26]
  PIN data_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.2691 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.896 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 30.0562 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 137.238 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 444.770000 550.160000 445.150000 ;
    END
  END data_rdata_i[25]
  PIN data_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.6023 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.536 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 33.2765 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 154.893 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.566667 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 447.210000 550.160000 447.590000 ;
    END
  END data_rdata_i[24]
  PIN data_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.6328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.512 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 59.4147 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 290.956 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.778944 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 449.650000 550.160000 450.030000 ;
    END
  END data_rdata_i[23]
  PIN data_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2106 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.2448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 81.776 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 52.4901 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 258.815 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.620214 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 452.090000 550.160000 452.470000 ;
    END
  END data_rdata_i[22]
  PIN data_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.3995 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.4 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 28.3822 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 130.556 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 453.920000 550.160000 454.300000 ;
    END
  END data_rdata_i[21]
  PIN data_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.2744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.792 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 41.536 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 196.771 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.461484 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 456.360000 550.160000 456.740000 ;
    END
  END data_rdata_i[20]
  PIN data_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 14.8048 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 56.4569 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.313033 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 458.800000 550.160000 459.180000 ;
    END
  END data_rdata_i[19]
  PIN data_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.816 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 35.5409 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 165.862 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.798786 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 461.240000 550.160000 461.620000 ;
    END
  END data_rdata_i[18]
  PIN data_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.496 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 26.1064 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 116.71 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.372198 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 463.070000 550.160000 463.450000 ;
    END
  END data_rdata_i[17]
  PIN data_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.1742 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 35.2093 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 163.415 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.944697 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 465.510000 550.160000 465.890000 ;
    END
  END data_rdata_i[16]
  PIN data_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9472 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 31.1673 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 142.288 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.461484 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 467.950000 550.160000 468.330000 ;
    END
  END data_rdata_i[15]
  PIN data_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.3946 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.9678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 117.632 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 44.8803 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 219.569 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.620214 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 470.390000 550.160000 470.770000 ;
    END
  END data_rdata_i[14]
  PIN data_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.2906 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 92.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.8088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 100.784 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 35.5877 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 170.364 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.515032 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 472.830000 550.160000 473.210000 ;
    END
  END data_rdata_i[13]
  PIN data_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0006 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 38.8215 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 207.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 68.0608 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 342.11 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 474.660000 550.160000 475.040000 ;
    END
  END data_rdata_i[12]
  PIN data_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.2246 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.2677 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 76.56 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 65.4472 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 321.377 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 477.100000 550.160000 477.480000 ;
    END
  END data_rdata_i[11]
  PIN data_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.32 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 28.6634 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 126.541 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.461484 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 479.540000 550.160000 479.920000 ;
    END
  END data_rdata_i[10]
  PIN data_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2044 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.752 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 15.2147 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 58.9259 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.372198 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 481.980000 550.160000 482.360000 ;
    END
  END data_rdata_i[9]
  PIN data_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.112 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 19.4692 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 79.7591 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.640055 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 483.810000 550.160000 484.190000 ;
    END
  END data_rdata_i[8]
  PIN data_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3586 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 30.5208 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 163.248 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 57.2311 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 283.802 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.693603 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 486.250000 550.160000 486.630000 ;
    END
  END data_rdata_i[7]
  PIN data_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 49.4394 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 229.336 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.640055 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 488.690000 550.160000 489.070000 ;
    END
  END data_rdata_i[6]
  PIN data_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6212 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.112 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 40.3055 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 185.711 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 491.130000 550.160000 491.510000 ;
    END
  END data_rdata_i[5]
  PIN data_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2456 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.4806 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 179.504 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 57.4641 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 288.252 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 492.960000 550.160000 493.340000 ;
    END
  END data_rdata_i[4]
  PIN data_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.224 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 32.0271 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 142.964 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.372198 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 495.400000 550.160000 495.780000 ;
    END
  END data_rdata_i[3]
  PIN data_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3476 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 38.5806 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 206.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 68.868 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 348.625 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 497.840000 550.160000 498.220000 ;
    END
  END data_rdata_i[2]
  PIN data_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.6252 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.8 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 44.4905 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 209.356 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.566667 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 500.280000 550.160000 500.660000 ;
    END
  END data_rdata_i[1]
  PIN data_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.2384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.4 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 45.9046 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 236.727 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.346263 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.3278 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.552 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 55.7143 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 289.675 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.884127 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 502.110000 550.160000 502.490000 ;
    END
  END data_rdata_i[0]
  PIN data_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 549.260000 504.550000 550.160000 504.930000 ;
    END
  END data_err_i
  PIN irq_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6255 LAYER met3  ;
    ANTENNAMAXAREACAR 18.5228 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 76.2446 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.412362 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 506.990000 550.160000 507.370000 ;
    END
  END irq_i
  PIN irq_id_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.624 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 27.3832 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 141.236 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 509.430000 550.160000 509.810000 ;
    END
  END irq_id_i[4]
  PIN irq_id_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.888 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 25.721 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 131.786 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 511.260000 550.160000 511.640000 ;
    END
  END irq_id_i[3]
  PIN irq_id_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.28 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 14.1505 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 69.8465 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 513.700000 550.160000 514.080000 ;
    END
  END irq_id_i[2]
  PIN irq_id_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9754 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.864 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 26.144 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 134.343 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 516.140000 550.160000 516.520000 ;
    END
  END irq_id_i[1]
  PIN irq_id_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 12.2337 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 57.7818 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 518.580000 550.160000 518.960000 ;
    END
  END irq_id_i[0]
  PIN irq_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 532.000000 550.160000 532.380000 ;
    END
  END irq_ack_o
  PIN irq_id_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 520.410000 550.160000 520.790000 ;
    END
  END irq_id_o[4]
  PIN irq_id_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.8944 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.432 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 522.850000 550.160000 523.230000 ;
    END
  END irq_id_o[3]
  PIN irq_id_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.4804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.224 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 525.290000 550.160000 525.670000 ;
    END
  END irq_id_o[2]
  PIN irq_id_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 527.730000 550.160000 528.110000 ;
    END
  END irq_id_o[1]
  PIN irq_id_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 529.560000 550.160000 529.940000 ;
    END
  END irq_id_o[0]
  PIN debug_req_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 40.9245 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 185.628 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.257516 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 534.440000 550.160000 534.820000 ;
    END
  END debug_req_i
  PIN fetch_enable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.196 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.648 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 36.6212 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 189.758 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 536.880000 550.160000 537.260000 ;
    END
  END fetch_enable_i
  PIN ext_perf_counters_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.2078 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 59.4314 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 327.321 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 538.710000 550.160000 539.090000 ;
    END
  END ext_perf_counters_i
  PIN eFPGA_operand_a_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4413 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.678 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.6318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 195.84 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 10.160000 0.000000 10.540000 0.900000 ;
    END
  END eFPGA_operand_a_o[31]
  PIN eFPGA_operand_a_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 12.920000 0.000000 13.300000 0.900000 ;
    END
  END eFPGA_operand_a_o[30]
  PIN eFPGA_operand_a_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4489 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.0835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.849 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 54.1278 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 289.152 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 16.140000 0.000000 16.520000 0.900000 ;
    END
  END eFPGA_operand_a_o[29]
  PIN eFPGA_operand_a_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 63.2538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 337.824 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 19.360000 0.000000 19.740000 0.900000 ;
    END
  END eFPGA_operand_a_o[28]
  PIN eFPGA_operand_a_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.8885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.2466 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 306.256 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 22.580000 0.000000 22.960000 0.900000 ;
    END
  END eFPGA_operand_a_o[27]
  PIN eFPGA_operand_a_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5567 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.6826 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 287.248 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 25.800000 0.000000 26.180000 0.900000 ;
    END
  END eFPGA_operand_a_o[26]
  PIN eFPGA_operand_a_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3921 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.9798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 277.696 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 29.020000 0.000000 29.400000 0.900000 ;
    END
  END eFPGA_operand_a_o[25]
  PIN eFPGA_operand_a_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0355 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.678 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 55.1388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 294.544 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 31.780000 0.000000 32.160000 0.900000 ;
    END
  END eFPGA_operand_a_o[24]
  PIN eFPGA_operand_a_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1267 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.3545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.526 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.9434 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 203.776 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 35.000000 0.000000 35.380000 0.900000 ;
    END
  END eFPGA_operand_a_o[23]
  PIN eFPGA_operand_a_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3749 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.5955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.223 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.9798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 309.696 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 38.220000 0.000000 38.600000 0.900000 ;
    END
  END eFPGA_operand_a_o[22]
  PIN eFPGA_operand_a_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7056 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.55131 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.9118 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0995286 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 41.440000 0.000000 41.820000 0.900000 ;
    END
  END eFPGA_operand_a_o[21]
  PIN eFPGA_operand_a_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.8238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 132.864 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 44.660000 0.000000 45.040000 0.900000 ;
    END
  END eFPGA_operand_a_o[20]
  PIN eFPGA_operand_a_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4413 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.9808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 112.368 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 47.880000 0.000000 48.260000 0.900000 ;
    END
  END eFPGA_operand_a_o[19]
  PIN eFPGA_operand_a_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4818 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.301 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 51.100000 0.000000 51.480000 0.900000 ;
    END
  END eFPGA_operand_a_o[18]
  PIN eFPGA_operand_a_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4818 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.301 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 53.860000 0.000000 54.240000 0.900000 ;
    END
  END eFPGA_operand_a_o[17]
  PIN eFPGA_operand_a_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.459 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 57.080000 0.000000 57.460000 0.900000 ;
    END
  END eFPGA_operand_a_o[16]
  PIN eFPGA_operand_a_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1641 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.666 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 121.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.2448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 65.776 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 60.300000 0.000000 60.680000 0.900000 ;
    END
  END eFPGA_operand_a_o[15]
  PIN eFPGA_operand_a_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.154 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 63.520000 0.000000 63.900000 0.900000 ;
    END
  END eFPGA_operand_a_o[14]
  PIN eFPGA_operand_a_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.488 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.5758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 78.208 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 66.740000 0.000000 67.120000 0.900000 ;
    END
  END eFPGA_operand_a_o[13]
  PIN eFPGA_operand_a_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9141 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.2915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 69.960000 0.000000 70.340000 0.900000 ;
    END
  END eFPGA_operand_a_o[12]
  PIN eFPGA_operand_a_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.992 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.734 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 73.180000 0.000000 73.560000 0.900000 ;
    END
  END eFPGA_operand_a_o[11]
  PIN eFPGA_operand_a_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8811 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.1968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 65.52 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 75.940000 0.000000 76.320000 0.900000 ;
    END
  END eFPGA_operand_a_o[10]
  PIN eFPGA_operand_a_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.7536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.542 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 79.160000 0.000000 79.540000 0.900000 ;
    END
  END eFPGA_operand_a_o[9]
  PIN eFPGA_operand_a_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.318 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.472 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 82.380000 0.000000 82.760000 0.900000 ;
    END
  END eFPGA_operand_a_o[8]
  PIN eFPGA_operand_a_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9562 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.555 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 85.600000 0.000000 85.980000 0.900000 ;
    END
  END eFPGA_operand_a_o[7]
  PIN eFPGA_operand_a_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7514 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.531 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 88.820000 0.000000 89.200000 0.900000 ;
    END
  END eFPGA_operand_a_o[6]
  PIN eFPGA_operand_a_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8683 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.6528 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 323.952 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 92.040000 0.000000 92.420000 0.900000 ;
    END
  END eFPGA_operand_a_o[5]
  PIN eFPGA_operand_a_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.5681 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.6795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.092 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.6048 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 323.696 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 94.800000 0.000000 95.180000 0.900000 ;
    END
  END eFPGA_operand_a_o[4]
  PIN eFPGA_operand_a_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6975 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 67.6938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 361.504 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 98.020000 0.000000 98.400000 0.900000 ;
    END
  END eFPGA_operand_a_o[3]
  PIN eFPGA_operand_a_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3749 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.5955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.8648 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 218.416 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 101.240000 0.000000 101.620000 0.900000 ;
    END
  END eFPGA_operand_a_o[2]
  PIN eFPGA_operand_a_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6593 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.1355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.1018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 267.68 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 104.460000 0.000000 104.840000 0.900000 ;
    END
  END eFPGA_operand_a_o[1]
  PIN eFPGA_operand_a_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6975 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.4538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 88.224 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 107.680000 0.000000 108.060000 0.900000 ;
    END
  END eFPGA_operand_a_o[0]
  PIN eFPGA_operand_b_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.6618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 276 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 110.900000 0.000000 111.280000 0.900000 ;
    END
  END eFPGA_operand_b_o[31]
  PIN eFPGA_operand_b_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8473 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 61.2726 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 327.728 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 114.120000 0.000000 114.500000 0.900000 ;
    END
  END eFPGA_operand_b_o[30]
  PIN eFPGA_operand_b_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.503 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 62.7378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 335.072 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 116.880000 0.000000 117.260000 0.900000 ;
    END
  END eFPGA_operand_b_o[29]
  PIN eFPGA_operand_b_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0371 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.0245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.9888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 229.744 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 120.100000 0.000000 120.480000 0.900000 ;
    END
  END eFPGA_operand_b_o[28]
  PIN eFPGA_operand_b_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.8405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.4438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 301.504 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 123.320000 0.000000 123.700000 0.900000 ;
    END
  END eFPGA_operand_b_o[27]
  PIN eFPGA_operand_b_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0615 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.438 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 62.2128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 332.272 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 126.540000 0.000000 126.920000 0.900000 ;
    END
  END eFPGA_operand_b_o[26]
  PIN eFPGA_operand_b_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1245 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.16 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.3718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 301.12 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 129.760000 0.000000 130.140000 0.900000 ;
    END
  END eFPGA_operand_b_o[25]
  PIN eFPGA_operand_b_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2781 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.2295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.2108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 278.928 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 132.980000 0.000000 133.360000 0.900000 ;
    END
  END eFPGA_operand_b_o[24]
  PIN eFPGA_operand_b_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0997 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.473 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 63.6528 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 339.952 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 136.200000 0.000000 136.580000 0.900000 ;
    END
  END eFPGA_operand_b_o[23]
  PIN eFPGA_operand_b_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.5457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.5675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.1978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 252.192 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 138.960000 0.000000 139.340000 0.900000 ;
    END
  END eFPGA_operand_b_o[22]
  PIN eFPGA_operand_b_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.7628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 153.872 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 142.180000 0.000000 142.560000 0.900000 ;
    END
  END eFPGA_operand_b_o[21]
  PIN eFPGA_operand_b_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4413 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.4558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 125.568 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 145.400000 0.000000 145.780000 0.900000 ;
    END
  END eFPGA_operand_b_o[20]
  PIN eFPGA_operand_b_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0925 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.3015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.332 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.2098 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 76.256 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 148.620000 0.000000 149.000000 0.900000 ;
    END
  END eFPGA_operand_b_o[19]
  PIN eFPGA_operand_b_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.1545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.16 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.6018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 115.68 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 151.840000 0.000000 152.220000 0.900000 ;
    END
  END eFPGA_operand_b_o[18]
  PIN eFPGA_operand_b_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.5668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 142.16 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 155.060000 0.000000 155.440000 0.900000 ;
    END
  END eFPGA_operand_b_o[17]
  PIN eFPGA_operand_b_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4366 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.075 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 158.280000 0.000000 158.660000 0.900000 ;
    END
  END eFPGA_operand_b_o[16]
  PIN eFPGA_operand_b_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 161.040000 0.000000 161.420000 0.900000 ;
    END
  END eFPGA_operand_b_o[15]
  PIN eFPGA_operand_b_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3174 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.361 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 164.260000 0.000000 164.640000 0.900000 ;
    END
  END eFPGA_operand_b_o[14]
  PIN eFPGA_operand_b_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4818 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.301 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 167.480000 0.000000 167.860000 0.900000 ;
    END
  END eFPGA_operand_b_o[13]
  PIN eFPGA_operand_b_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4342 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.063 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 170.700000 0.000000 171.080000 0.900000 ;
    END
  END eFPGA_operand_b_o[12]
  PIN eFPGA_operand_b_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0997 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.9898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 80.416 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 173.920000 0.000000 174.300000 0.900000 ;
    END
  END eFPGA_operand_b_o[11]
  PIN eFPGA_operand_b_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.0634 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.091 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 177.140000 0.000000 177.520000 0.900000 ;
    END
  END eFPGA_operand_b_o[10]
  PIN eFPGA_operand_b_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.8608 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.078 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 179.900000 0.000000 180.280000 0.900000 ;
    END
  END eFPGA_operand_b_o[9]
  PIN eFPGA_operand_b_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.337 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.577 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 183.120000 0.000000 183.500000 0.900000 ;
    END
  END eFPGA_operand_b_o[8]
  PIN eFPGA_operand_b_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.437 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 186.340000 0.000000 186.720000 0.900000 ;
    END
  END eFPGA_operand_b_o[7]
  PIN eFPGA_operand_b_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2533 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.1055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.5228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 216.592 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 189.560000 0.000000 189.940000 0.900000 ;
    END
  END eFPGA_operand_b_o[6]
  PIN eFPGA_operand_b_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1851 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.825 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.9946 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 208.912 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 192.780000 0.000000 193.160000 0.900000 ;
    END
  END eFPGA_operand_b_o[5]
  PIN eFPGA_operand_b_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0997 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.9018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 245.28 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 196.000000 0.000000 196.380000 0.900000 ;
    END
  END eFPGA_operand_b_o[4]
  PIN eFPGA_operand_b_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6121 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.5618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 232.8 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 199.220000 0.000000 199.600000 0.900000 ;
    END
  END eFPGA_operand_b_o[3]
  PIN eFPGA_operand_b_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.2938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 236.704 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 201.980000 0.000000 202.360000 0.900000 ;
    END
  END eFPGA_operand_b_o[2]
  PIN eFPGA_operand_b_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6975 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.1888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 300.144 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 205.200000 0.000000 205.580000 0.900000 ;
    END
  END eFPGA_operand_b_o[1]
  PIN eFPGA_operand_b_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6121 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.9718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 192.32 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 208.420000 0.000000 208.800000 0.900000 ;
    END
  END eFPGA_operand_b_o[0]
  PIN eFPGA_result_a_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1851 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 149.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 14.6604 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 74.2263 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 211.640000 0.000000 212.020000 0.900000 ;
    END
  END eFPGA_result_a_i[31]
  PIN eFPGA_result_a_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.863 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 10.3648 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 45.8323 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 214.860000 0.000000 215.240000 0.900000 ;
    END
  END eFPGA_result_a_i[30]
  PIN eFPGA_result_a_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6202 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.875 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.24465 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.1131 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 218.080000 0.000000 218.460000 0.900000 ;
    END
  END eFPGA_result_a_i[29]
  PIN eFPGA_result_a_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1176 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.362 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 6.21394 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.9596 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 221.300000 0.000000 221.680000 0.900000 ;
    END
  END eFPGA_result_a_i[28]
  PIN eFPGA_result_a_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.632 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 4.43434 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 16.6162 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 224.060000 0.000000 224.440000 0.900000 ;
    END
  END eFPGA_result_a_i[27]
  PIN eFPGA_result_a_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9128 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.338 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.42687 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.0242 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 227.280000 0.000000 227.660000 0.900000 ;
    END
  END eFPGA_result_a_i[26]
  PIN eFPGA_result_a_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0624 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.968 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 10.0313 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.5697 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 230.500000 0.000000 230.880000 0.900000 ;
    END
  END eFPGA_result_a_i[25]
  PIN eFPGA_result_a_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6563 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.336 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 16.9758 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 87.3273 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 233.720000 0.000000 234.100000 0.900000 ;
    END
  END eFPGA_result_a_i[24]
  PIN eFPGA_result_a_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1489 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.5735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 57.5438 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 301.392 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 236.940000 0.000000 237.320000 0.900000 ;
    END
  END eFPGA_result_a_i[23]
  PIN eFPGA_result_a_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2702 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.125 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 7.70909 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.5535 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 240.160000 0.000000 240.540000 0.900000 ;
    END
  END eFPGA_result_a_i[22]
  PIN eFPGA_result_a_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7619 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.308 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 156.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 11.5 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 60.5697 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 242.920000 0.000000 243.300000 0.900000 ;
    END
  END eFPGA_result_a_i[21]
  PIN eFPGA_result_a_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3233 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.1034 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 55.296 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 44.3921 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 237.895 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 246.140000 0.000000 246.520000 0.900000 ;
    END
  END eFPGA_result_a_i[20]
  PIN eFPGA_result_a_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9472 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.618 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.50949 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 42.1556 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 249.360000 0.000000 249.740000 0.900000 ;
    END
  END eFPGA_result_a_i[19]
  PIN eFPGA_result_a_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3315 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.3785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 18.7137 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 101.939 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 252.580000 0.000000 252.960000 0.900000 ;
    END
  END eFPGA_result_a_i[18]
  PIN eFPGA_result_a_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6986 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.267 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.85576 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.2869 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 255.800000 0.000000 256.180000 0.900000 ;
    END
  END eFPGA_result_a_i[17]
  PIN eFPGA_result_a_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1274 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.411 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 6.50707 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.5434 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 259.020000 0.000000 259.400000 0.900000 ;
    END
  END eFPGA_result_a_i[16]
  PIN eFPGA_result_a_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6962 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.137 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 18.2917 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 84.9899 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 262.240000 0.000000 262.620000 0.900000 ;
    END
  END eFPGA_result_a_i[15]
  PIN eFPGA_result_a_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.6565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.798 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.056 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 17.8061 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 90.1657 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 265.000000 0.000000 265.380000 0.900000 ;
    END
  END eFPGA_result_a_i[14]
  PIN eFPGA_result_a_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8044 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.904 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.93253 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.2707 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 268.220000 0.000000 268.600000 0.900000 ;
    END
  END eFPGA_result_a_i[13]
  PIN eFPGA_result_a_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.991 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 117.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 28.6069 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 152.376 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 271.440000 0.000000 271.820000 0.900000 ;
    END
  END eFPGA_result_a_i[12]
  PIN eFPGA_result_a_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0696 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.122 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 10.0604 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.1919 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 274.660000 0.000000 275.040000 0.900000 ;
    END
  END eFPGA_result_a_i[11]
  PIN eFPGA_result_a_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.9658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.288 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 86.7665 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 453.683 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 277.880000 0.000000 278.260000 0.900000 ;
    END
  END eFPGA_result_a_i[10]
  PIN eFPGA_result_a_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5972 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.868 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.65535 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 42.7212 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 281.100000 0.000000 281.480000 0.900000 ;
    END
  END eFPGA_result_a_i[9]
  PIN eFPGA_result_a_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.889 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.219 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 11.0945 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 49.4808 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 284.320000 0.000000 284.700000 0.900000 ;
    END
  END eFPGA_result_a_i[8]
  PIN eFPGA_result_a_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9803 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.6225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.652 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 147.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 22.4964 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 114.255 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 287.080000 0.000000 287.460000 0.900000 ;
    END
  END eFPGA_result_a_i[7]
  PIN eFPGA_result_a_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7829 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.5972 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.4 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 25.564 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 138.733 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 290.300000 0.000000 290.680000 0.900000 ;
    END
  END eFPGA_result_a_i[6]
  PIN eFPGA_result_a_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.863 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 10.3139 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 45.5778 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 293.520000 0.000000 293.900000 0.900000 ;
    END
  END eFPGA_result_a_i[5]
  PIN eFPGA_result_a_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.001 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.779 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.78323 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 42.8061 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 296.740000 0.000000 297.120000 0.900000 ;
    END
  END eFPGA_result_a_i[4]
  PIN eFPGA_result_a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.651 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.029 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.88283 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.4222 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 299.960000 0.000000 300.340000 0.900000 ;
    END
  END eFPGA_result_a_i[3]
  PIN eFPGA_result_a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6412 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.98 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.32949 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.5374 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 303.180000 0.000000 303.560000 0.900000 ;
    END
  END eFPGA_result_a_i[2]
  PIN eFPGA_result_a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.671 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 94.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 16.8123 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 88.497 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 306.400000 0.000000 306.780000 0.900000 ;
    END
  END eFPGA_result_a_i[1]
  PIN eFPGA_result_a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3067 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.3725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 35.971 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 192.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.4868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.4 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 35.3368 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 184.933 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 309.160000 0.000000 309.540000 0.900000 ;
    END
  END eFPGA_result_a_i[0]
  PIN eFPGA_result_b_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1482 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.633 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 27.7484 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 120.107 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 312.380000 0.000000 312.760000 0.900000 ;
    END
  END eFPGA_result_b_i[31]
  PIN eFPGA_result_b_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7504 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.526 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 23.8357 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 99.6071 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 315.600000 0.000000 315.980000 0.900000 ;
    END
  END eFPGA_result_b_i[30]
  PIN eFPGA_result_b_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3246 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.515 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 32.3484 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 143.107 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 318.820000 0.000000 319.200000 0.900000 ;
    END
  END eFPGA_result_b_i[29]
  PIN eFPGA_result_b_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6578 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.181 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 26.5524 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 114.663 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 322.040000 0.000000 322.420000 0.900000 ;
    END
  END eFPGA_result_b_i[28]
  PIN eFPGA_result_b_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.643 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 27.6817 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 119.774 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 325.260000 0.000000 325.640000 0.900000 ;
    END
  END eFPGA_result_b_i[27]
  PIN eFPGA_result_b_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2602 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.193 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 25.704 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 109.885 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 328.020000 0.000000 328.400000 0.900000 ;
    END
  END eFPGA_result_b_i[26]
  PIN eFPGA_result_b_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0694 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.239 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 30.2151 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 132.44 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 331.240000 0.000000 331.620000 0.900000 ;
    END
  END eFPGA_result_b_i[25]
  PIN eFPGA_result_b_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.501 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.397 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 25.3079 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 108.44 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 334.460000 0.000000 334.840000 0.900000 ;
    END
  END eFPGA_result_b_i[24]
  PIN eFPGA_result_b_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6578 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.181 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 27.4595 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 118.663 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 337.680000 0.000000 338.060000 0.900000 ;
    END
  END eFPGA_result_b_i[23]
  PIN eFPGA_result_b_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.859 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 26.0413 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 112.107 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 340.900000 0.000000 341.280000 0.900000 ;
    END
  END eFPGA_result_b_i[22]
  PIN eFPGA_result_b_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4842 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.313 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 27.6151 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 119.44 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 344.120000 0.000000 344.500000 0.900000 ;
    END
  END eFPGA_result_b_i[21]
  PIN eFPGA_result_b_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9742 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.763 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 35.3262 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 157.996 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 347.340000 0.000000 347.720000 0.900000 ;
    END
  END eFPGA_result_b_i[20]
  PIN eFPGA_result_b_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.477 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 31.6151 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 139.44 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 350.100000 0.000000 350.480000 0.900000 ;
    END
  END eFPGA_result_b_i[19]
  PIN eFPGA_result_b_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2434 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.109 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 23.2635 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 98.2183 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 353.320000 0.000000 353.700000 0.900000 ;
    END
  END eFPGA_result_b_i[18]
  PIN eFPGA_result_b_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0558 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.171 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 22.1706 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 92.2183 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 356.540000 0.000000 356.920000 0.900000 ;
    END
  END eFPGA_result_b_i[17]
  PIN eFPGA_result_b_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4366 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.075 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 24.7968 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 105.885 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 359.760000 0.000000 360.140000 0.900000 ;
    END
  END eFPGA_result_b_i[16]
  PIN eFPGA_result_b_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3722 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.753 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 24.6817 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 104.774 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 362.980000 0.000000 363.360000 0.900000 ;
    END
  END eFPGA_result_b_i[15]
  PIN eFPGA_result_b_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7674 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.729 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 21.9262 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 90.996 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 366.200000 0.000000 366.580000 0.900000 ;
    END
  END eFPGA_result_b_i[14]
  PIN eFPGA_result_b_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.277 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.277 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 25.704 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 109.885 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 369.420000 0.000000 369.800000 0.900000 ;
    END
  END eFPGA_result_b_i[13]
  PIN eFPGA_result_b_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.431 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 24.6817 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 104.774 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 372.180000 0.000000 372.560000 0.900000 ;
    END
  END eFPGA_result_b_i[12]
  PIN eFPGA_result_b_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.431 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 25.704 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 109.885 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 375.400000 0.000000 375.780000 0.900000 ;
    END
  END eFPGA_result_b_i[11]
  PIN eFPGA_result_b_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.859 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 26.0413 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 112.107 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 378.620000 0.000000 379.000000 0.900000 ;
    END
  END eFPGA_result_b_i[10]
  PIN eFPGA_result_b_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3722 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.753 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 24.6817 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 104.774 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 381.840000 0.000000 382.220000 0.900000 ;
    END
  END eFPGA_result_b_i[9]
  PIN eFPGA_result_b_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.859 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 29.404 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 128.385 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 385.060000 0.000000 385.440000 0.900000 ;
    END
  END eFPGA_result_b_i[8]
  PIN eFPGA_result_b_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5773 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.7785 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 26.3095 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 112.913 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 388.280000 0.000000 388.660000 0.900000 ;
    END
  END eFPGA_result_b_i[7]
  PIN eFPGA_result_b_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7222 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.503 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 27.0635 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 117.218 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 391.040000 0.000000 391.420000 0.900000 ;
    END
  END eFPGA_result_b_i[6]
  PIN eFPGA_result_b_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.085 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 33.2817 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 147.774 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 394.260000 0.000000 394.640000 0.900000 ;
    END
  END eFPGA_result_b_i[5]
  PIN eFPGA_result_b_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7222 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.503 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 27.0635 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 117.218 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 397.480000 0.000000 397.860000 0.900000 ;
    END
  END eFPGA_result_b_i[4]
  PIN eFPGA_result_b_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.441 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 32.804 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 145.385 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 400.700000 0.000000 401.080000 0.900000 ;
    END
  END eFPGA_result_b_i[3]
  PIN eFPGA_result_b_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.277 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.277 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 28.2595 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 122.663 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 403.920000 0.000000 404.300000 0.900000 ;
    END
  END eFPGA_result_b_i[2]
  PIN eFPGA_result_b_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.005 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.917 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 36.4929 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 163.829 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 407.140000 0.000000 407.520000 0.900000 ;
    END
  END eFPGA_result_b_i[1]
  PIN eFPGA_result_b_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9914 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.849 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 30.1151 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 131.94 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 410.360000 0.000000 410.740000 0.900000 ;
    END
  END eFPGA_result_b_i[0]
  PIN eFPGA_result_c_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3993 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.937 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 10.3861 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 56.5212 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 413.120000 0.000000 413.500000 0.900000 ;
    END
  END eFPGA_result_c_i[31]
  PIN eFPGA_result_c_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2181 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.8115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.1588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.984 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 48.2446 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 256.21 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 416.340000 0.000000 416.720000 0.900000 ;
    END
  END eFPGA_result_c_i[30]
  PIN eFPGA_result_c_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.108 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 3.43535 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.4485 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 419.560000 0.000000 419.940000 0.900000 ;
    END
  END eFPGA_result_c_i[29]
  PIN eFPGA_result_c_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0318 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.933 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 16.4741 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 79.9333 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 422.780000 0.000000 423.160000 0.900000 ;
    END
  END eFPGA_result_c_i[28]
  PIN eFPGA_result_c_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9846 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.697 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 4.80667 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.8687 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 426.000000 0.000000 426.380000 0.900000 ;
    END
  END eFPGA_result_c_i[27]
  PIN eFPGA_result_c_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.2828 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 49.0552 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 259.083 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 429.220000 0.000000 429.600000 0.900000 ;
    END
  END eFPGA_result_c_i[26]
  PIN eFPGA_result_c_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.3865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.202 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 161.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.816 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 20.9509 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 112.299 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 432.440000 0.000000 432.820000 0.900000 ;
    END
  END eFPGA_result_c_i[25]
  PIN eFPGA_result_c_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9846 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.697 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 5.21758 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.6505 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 435.200000 0.000000 435.580000 0.900000 ;
    END
  END eFPGA_result_c_i[24]
  PIN eFPGA_result_c_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9842 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.695 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.56747 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 45.4 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 438.420000 0.000000 438.800000 0.900000 ;
    END
  END eFPGA_result_c_i[23]
  PIN eFPGA_result_c_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5553 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.6155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.187 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 145.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 29.561 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 157.616 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 441.640000 0.000000 442.020000 0.900000 ;
    END
  END eFPGA_result_c_i[22]
  PIN eFPGA_result_c_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4481 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 6.57677 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 34.901 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 444.860000 0.000000 445.240000 0.900000 ;
    END
  END eFPGA_result_c_i[21]
  PIN eFPGA_result_c_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.435 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 7.82727 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 36.9717 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 448.080000 0.000000 448.460000 0.900000 ;
    END
  END eFPGA_result_c_i[20]
  PIN eFPGA_result_c_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3807 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.337 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 98.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 14.6208 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 78.6182 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 451.300000 0.000000 451.680000 0.900000 ;
    END
  END eFPGA_result_c_i[19]
  PIN eFPGA_result_c_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7798 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.673 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.22121 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.6687 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 454.520000 0.000000 454.900000 0.900000 ;
    END
  END eFPGA_result_c_i[18]
  PIN eFPGA_result_c_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8894 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.221 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 4.42202 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.9455 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 457.280000 0.000000 457.660000 0.900000 ;
    END
  END eFPGA_result_c_i[17]
  PIN eFPGA_result_c_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9912 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.73 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.28465 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.9859 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 460.500000 0.000000 460.880000 0.900000 ;
    END
  END eFPGA_result_c_i[16]
  PIN eFPGA_result_c_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.113 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.339 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.82768 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.701 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 463.720000 0.000000 464.100000 0.900000 ;
    END
  END eFPGA_result_c_i[15]
  PIN eFPGA_result_c_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8418 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.983 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 4.2297 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.9838 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 466.940000 0.000000 467.320000 0.900000 ;
    END
  END eFPGA_result_c_i[14]
  PIN eFPGA_result_c_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0794 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.171 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 10.4046 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 49.5859 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 470.160000 0.000000 470.540000 0.900000 ;
    END
  END eFPGA_result_c_i[13]
  PIN eFPGA_result_c_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.525 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 120.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 13.5335 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 73.4788 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 473.380000 0.000000 473.760000 0.900000 ;
    END
  END eFPGA_result_c_i[12]
  PIN eFPGA_result_c_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6975 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 13.6475 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 79.6242 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 476.140000 0.000000 476.520000 0.900000 ;
    END
  END eFPGA_result_c_i[11]
  PIN eFPGA_result_c_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3559 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.361 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 162.392 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 9.89879 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 54.0444 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 479.360000 0.000000 479.740000 0.900000 ;
    END
  END eFPGA_result_c_i[10]
  PIN eFPGA_result_c_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.963 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.471 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.7598 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.1576 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 482.580000 0.000000 482.960000 0.900000 ;
    END
  END eFPGA_result_c_i[9]
  PIN eFPGA_result_c_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3251 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.3365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.677 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.8204 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.12 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 46.3376 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 252.186 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 485.800000 0.000000 486.180000 0.900000 ;
    END
  END eFPGA_result_c_i[8]
  PIN eFPGA_result_c_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5558 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.553 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.80949 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.6101 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 489.020000 0.000000 489.400000 0.900000 ;
    END
  END eFPGA_result_c_i[7]
  PIN eFPGA_result_c_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5267 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.339 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 119.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 15.382 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 80.105 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 492.240000 0.000000 492.620000 0.900000 ;
    END
  END eFPGA_result_c_i[6]
  PIN eFPGA_result_c_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2533 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.1055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 13.6232 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 79.4101 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 495.460000 0.000000 495.840000 0.900000 ;
    END
  END eFPGA_result_c_i[5]
  PIN eFPGA_result_c_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3559 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.7146 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.752 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 21.8257 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 117.871 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 498.220000 0.000000 498.600000 0.900000 ;
    END
  END eFPGA_result_c_i[4]
  PIN eFPGA_result_c_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4172 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.86 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 6.55455 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.6081 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 501.440000 0.000000 501.820000 0.900000 ;
    END
  END eFPGA_result_c_i[3]
  PIN eFPGA_result_c_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0798 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.173 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 5.19131 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.7919 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 504.660000 0.000000 505.040000 0.900000 ;
    END
  END eFPGA_result_c_i[2]
  PIN eFPGA_result_c_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.978 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.772 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.8204 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 42.3737 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 507.880000 0.000000 508.260000 0.900000 ;
    END
  END eFPGA_result_c_i[1]
  PIN eFPGA_result_c_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3559 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 15.3408 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 83.1515 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 511.100000 0.000000 511.480000 0.900000 ;
    END
  END eFPGA_result_c_i[0]
  PIN eFPGA_write_strobe_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0318 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.933 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 514.320000 0.000000 514.700000 0.900000 ;
    END
  END eFPGA_write_strobe_o
  PIN eFPGA_fpga_done_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.91 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.324 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 14.6043 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 55.3104 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.265597 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 517.540000 0.000000 517.920000 0.900000 ;
    END
  END eFPGA_fpga_done_i
  PIN eFPGA_en_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7672 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.61 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 520.300000 0.000000 520.680000 0.900000 ;
    END
  END eFPGA_en_o
  PIN eFPGA_operator_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1816 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.682 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 523.520000 0.000000 523.900000 0.900000 ;
    END
  END eFPGA_operator_o[1]
  PIN eFPGA_operator_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1851 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 28.1748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 150.736 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 526.740000 0.000000 527.120000 0.900000 ;
    END
  END eFPGA_operator_o[0]
  PIN eFPGA_delay_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.4318 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.933 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 529.960000 0.000000 530.340000 0.900000 ;
    END
  END eFPGA_delay_o[3]
  PIN eFPGA_delay_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.599 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 533.180000 0.000000 533.560000 0.900000 ;
    END
  END eFPGA_delay_o[2]
  PIN eFPGA_delay_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.921 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 536.400000 0.000000 536.780000 0.900000 ;
    END
  END eFPGA_delay_o[1]
  PIN eFPGA_delay_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.7598 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.856 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 539.160000 0.000000 539.540000 0.900000 ;
    END
  END eFPGA_delay_o[0]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 548.160000 541.160000 550.160000 543.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 541.160000 2.000000 543.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 548.160000 5.430000 550.160000 7.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 5.430000 2.000000 7.430000 ;
    END
    PORT
      LAYER met4 ;
        RECT 542.600000 547.780000 544.600000 549.780000 ;
    END
    PORT
      LAYER met4 ;
        RECT 542.600000 0.000000 544.600000 2.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 5.560000 547.780000 7.560000 549.780000 ;
    END
    PORT
      LAYER met4 ;
        RECT 5.560000 0.000000 7.560000 2.000000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 5.430000 550.160000 7.430000 ;
        RECT 0.000000 541.160000 550.160000 543.160000 ;
        RECT 5.560000 9.620000 7.560000 10.100000 ;
        RECT 5.560000 15.060000 7.560000 15.540000 ;
        RECT 12.120000 9.620000 13.320000 10.100000 ;
        RECT 12.120000 15.060000 13.320000 15.540000 ;
        RECT 5.560000 20.500000 7.560000 20.980000 ;
        RECT 12.120000 20.500000 13.320000 20.980000 ;
        RECT 5.560000 25.940000 7.560000 26.420000 ;
        RECT 5.560000 31.380000 7.560000 31.860000 ;
        RECT 12.120000 31.380000 13.320000 31.860000 ;
        RECT 12.120000 25.940000 13.320000 26.420000 ;
        RECT 57.120000 31.380000 58.320000 31.860000 ;
        RECT 57.120000 25.940000 58.320000 26.420000 ;
        RECT 57.120000 20.500000 58.320000 20.980000 ;
        RECT 57.120000 15.060000 58.320000 15.540000 ;
        RECT 57.120000 9.620000 58.320000 10.100000 ;
        RECT 5.560000 36.820000 7.560000 37.300000 ;
        RECT 5.560000 42.260000 7.560000 42.740000 ;
        RECT 12.120000 42.260000 13.320000 42.740000 ;
        RECT 12.120000 36.820000 13.320000 37.300000 ;
        RECT 5.560000 47.700000 7.560000 48.180000 ;
        RECT 12.120000 47.700000 13.320000 48.180000 ;
        RECT 5.560000 53.140000 7.560000 53.620000 ;
        RECT 5.560000 58.580000 7.560000 59.060000 ;
        RECT 12.120000 58.580000 13.320000 59.060000 ;
        RECT 12.120000 53.140000 13.320000 53.620000 ;
        RECT 5.560000 64.020000 7.560000 64.500000 ;
        RECT 12.120000 64.020000 13.320000 64.500000 ;
        RECT 57.120000 47.700000 58.320000 48.180000 ;
        RECT 57.120000 42.260000 58.320000 42.740000 ;
        RECT 57.120000 36.820000 58.320000 37.300000 ;
        RECT 57.120000 58.580000 58.320000 59.060000 ;
        RECT 57.120000 53.140000 58.320000 53.620000 ;
        RECT 57.120000 64.020000 58.320000 64.500000 ;
        RECT 102.120000 9.620000 103.320000 10.100000 ;
        RECT 102.120000 15.060000 103.320000 15.540000 ;
        RECT 102.120000 20.500000 103.320000 20.980000 ;
        RECT 102.120000 25.940000 103.320000 26.420000 ;
        RECT 102.120000 31.380000 103.320000 31.860000 ;
        RECT 102.120000 64.020000 103.320000 64.500000 ;
        RECT 102.120000 36.820000 103.320000 37.300000 ;
        RECT 102.120000 42.260000 103.320000 42.740000 ;
        RECT 102.120000 47.700000 103.320000 48.180000 ;
        RECT 102.120000 53.140000 103.320000 53.620000 ;
        RECT 102.120000 58.580000 103.320000 59.060000 ;
        RECT 5.560000 69.460000 7.560000 69.940000 ;
        RECT 5.560000 74.900000 7.560000 75.380000 ;
        RECT 12.120000 74.900000 13.320000 75.380000 ;
        RECT 12.120000 69.460000 13.320000 69.940000 ;
        RECT 5.560000 80.340000 7.560000 80.820000 ;
        RECT 12.120000 80.340000 13.320000 80.820000 ;
        RECT 5.560000 85.780000 7.560000 86.260000 ;
        RECT 12.120000 85.780000 13.320000 86.260000 ;
        RECT 12.120000 91.220000 13.320000 91.700000 ;
        RECT 5.560000 91.220000 7.560000 91.700000 ;
        RECT 5.560000 96.660000 7.560000 97.140000 ;
        RECT 5.560000 102.100000 7.560000 102.580000 ;
        RECT 12.120000 96.660000 13.320000 97.140000 ;
        RECT 12.120000 102.100000 13.320000 102.580000 ;
        RECT 57.120000 80.340000 58.320000 80.820000 ;
        RECT 57.120000 74.900000 58.320000 75.380000 ;
        RECT 57.120000 69.460000 58.320000 69.940000 ;
        RECT 57.120000 85.780000 58.320000 86.260000 ;
        RECT 57.120000 91.220000 58.320000 91.700000 ;
        RECT 57.120000 96.660000 58.320000 97.140000 ;
        RECT 57.120000 102.100000 58.320000 102.580000 ;
        RECT 5.560000 107.540000 7.560000 108.020000 ;
        RECT 12.120000 107.540000 13.320000 108.020000 ;
        RECT 5.560000 112.980000 7.560000 113.460000 ;
        RECT 5.560000 118.420000 7.560000 118.900000 ;
        RECT 12.120000 118.420000 13.320000 118.900000 ;
        RECT 12.120000 112.980000 13.320000 113.460000 ;
        RECT 5.560000 123.860000 7.560000 124.340000 ;
        RECT 12.120000 123.860000 13.320000 124.340000 ;
        RECT 5.560000 129.300000 7.560000 129.780000 ;
        RECT 5.560000 134.740000 7.560000 135.220000 ;
        RECT 12.120000 129.300000 13.320000 129.780000 ;
        RECT 12.120000 134.740000 13.320000 135.220000 ;
        RECT 57.120000 118.420000 58.320000 118.900000 ;
        RECT 57.120000 112.980000 58.320000 113.460000 ;
        RECT 57.120000 107.540000 58.320000 108.020000 ;
        RECT 57.120000 129.300000 58.320000 129.780000 ;
        RECT 57.120000 123.860000 58.320000 124.340000 ;
        RECT 57.120000 134.740000 58.320000 135.220000 ;
        RECT 102.120000 80.340000 103.320000 80.820000 ;
        RECT 102.120000 74.900000 103.320000 75.380000 ;
        RECT 102.120000 69.460000 103.320000 69.940000 ;
        RECT 102.120000 85.780000 103.320000 86.260000 ;
        RECT 102.120000 91.220000 103.320000 91.700000 ;
        RECT 102.120000 96.660000 103.320000 97.140000 ;
        RECT 102.120000 102.100000 103.320000 102.580000 ;
        RECT 102.120000 134.740000 103.320000 135.220000 ;
        RECT 102.120000 129.300000 103.320000 129.780000 ;
        RECT 102.120000 123.860000 103.320000 124.340000 ;
        RECT 102.120000 107.540000 103.320000 108.020000 ;
        RECT 102.120000 112.980000 103.320000 113.460000 ;
        RECT 102.120000 118.420000 103.320000 118.900000 ;
        RECT 147.120000 31.380000 148.320000 31.860000 ;
        RECT 147.120000 25.940000 148.320000 26.420000 ;
        RECT 147.120000 20.500000 148.320000 20.980000 ;
        RECT 147.120000 15.060000 148.320000 15.540000 ;
        RECT 147.120000 9.620000 148.320000 10.100000 ;
        RECT 192.120000 31.380000 193.320000 31.860000 ;
        RECT 192.120000 25.940000 193.320000 26.420000 ;
        RECT 192.120000 15.060000 193.320000 15.540000 ;
        RECT 192.120000 9.620000 193.320000 10.100000 ;
        RECT 192.120000 20.500000 193.320000 20.980000 ;
        RECT 147.120000 47.700000 148.320000 48.180000 ;
        RECT 147.120000 42.260000 148.320000 42.740000 ;
        RECT 147.120000 36.820000 148.320000 37.300000 ;
        RECT 147.120000 58.580000 148.320000 59.060000 ;
        RECT 147.120000 53.140000 148.320000 53.620000 ;
        RECT 147.120000 64.020000 148.320000 64.500000 ;
        RECT 192.120000 47.700000 193.320000 48.180000 ;
        RECT 192.120000 42.260000 193.320000 42.740000 ;
        RECT 192.120000 36.820000 193.320000 37.300000 ;
        RECT 192.120000 58.580000 193.320000 59.060000 ;
        RECT 192.120000 53.140000 193.320000 53.620000 ;
        RECT 192.120000 64.020000 193.320000 64.500000 ;
        RECT 237.120000 9.620000 238.320000 10.100000 ;
        RECT 237.120000 15.060000 238.320000 15.540000 ;
        RECT 237.120000 20.500000 238.320000 20.980000 ;
        RECT 237.120000 25.940000 238.320000 26.420000 ;
        RECT 237.120000 31.380000 238.320000 31.860000 ;
        RECT 237.120000 36.820000 238.320000 37.300000 ;
        RECT 237.120000 42.260000 238.320000 42.740000 ;
        RECT 237.120000 47.700000 238.320000 48.180000 ;
        RECT 237.120000 64.020000 238.320000 64.500000 ;
        RECT 237.120000 53.140000 238.320000 53.620000 ;
        RECT 237.120000 58.580000 238.320000 59.060000 ;
        RECT 147.120000 80.340000 148.320000 80.820000 ;
        RECT 147.120000 74.900000 148.320000 75.380000 ;
        RECT 147.120000 69.460000 148.320000 69.940000 ;
        RECT 147.120000 96.660000 148.320000 97.140000 ;
        RECT 147.120000 85.780000 148.320000 86.260000 ;
        RECT 147.120000 91.220000 148.320000 91.700000 ;
        RECT 147.120000 102.100000 148.320000 102.580000 ;
        RECT 192.120000 80.340000 193.320000 80.820000 ;
        RECT 192.120000 74.900000 193.320000 75.380000 ;
        RECT 192.120000 69.460000 193.320000 69.940000 ;
        RECT 192.120000 85.780000 193.320000 86.260000 ;
        RECT 192.120000 91.220000 193.320000 91.700000 ;
        RECT 192.120000 96.660000 193.320000 97.140000 ;
        RECT 192.120000 102.100000 193.320000 102.580000 ;
        RECT 147.120000 118.420000 148.320000 118.900000 ;
        RECT 147.120000 112.980000 148.320000 113.460000 ;
        RECT 147.120000 107.540000 148.320000 108.020000 ;
        RECT 147.120000 129.300000 148.320000 129.780000 ;
        RECT 147.120000 123.860000 148.320000 124.340000 ;
        RECT 147.120000 134.740000 148.320000 135.220000 ;
        RECT 192.120000 118.420000 193.320000 118.900000 ;
        RECT 192.120000 112.980000 193.320000 113.460000 ;
        RECT 192.120000 107.540000 193.320000 108.020000 ;
        RECT 192.120000 129.300000 193.320000 129.780000 ;
        RECT 192.120000 123.860000 193.320000 124.340000 ;
        RECT 192.120000 134.740000 193.320000 135.220000 ;
        RECT 237.120000 80.340000 238.320000 80.820000 ;
        RECT 237.120000 74.900000 238.320000 75.380000 ;
        RECT 237.120000 69.460000 238.320000 69.940000 ;
        RECT 237.120000 85.780000 238.320000 86.260000 ;
        RECT 237.120000 91.220000 238.320000 91.700000 ;
        RECT 237.120000 96.660000 238.320000 97.140000 ;
        RECT 237.120000 102.100000 238.320000 102.580000 ;
        RECT 237.120000 107.540000 238.320000 108.020000 ;
        RECT 237.120000 112.980000 238.320000 113.460000 ;
        RECT 237.120000 118.420000 238.320000 118.900000 ;
        RECT 237.120000 134.740000 238.320000 135.220000 ;
        RECT 237.120000 129.300000 238.320000 129.780000 ;
        RECT 237.120000 123.860000 238.320000 124.340000 ;
        RECT 12.120000 145.620000 13.320000 146.100000 ;
        RECT 5.560000 145.620000 7.560000 146.100000 ;
        RECT 12.120000 140.180000 13.320000 140.660000 ;
        RECT 5.560000 140.180000 7.560000 140.660000 ;
        RECT 5.560000 151.060000 7.560000 151.540000 ;
        RECT 12.120000 151.060000 13.320000 151.540000 ;
        RECT 5.560000 156.500000 7.560000 156.980000 ;
        RECT 5.560000 161.940000 7.560000 162.420000 ;
        RECT 12.120000 156.500000 13.320000 156.980000 ;
        RECT 12.120000 161.940000 13.320000 162.420000 ;
        RECT 5.560000 167.380000 7.560000 167.860000 ;
        RECT 12.120000 167.380000 13.320000 167.860000 ;
        RECT 57.120000 145.620000 58.320000 146.100000 ;
        RECT 57.120000 140.180000 58.320000 140.660000 ;
        RECT 57.120000 151.060000 58.320000 151.540000 ;
        RECT 57.120000 156.500000 58.320000 156.980000 ;
        RECT 57.120000 161.940000 58.320000 162.420000 ;
        RECT 57.120000 167.380000 58.320000 167.860000 ;
        RECT 5.560000 172.820000 7.560000 173.300000 ;
        RECT 5.560000 178.260000 7.560000 178.740000 ;
        RECT 12.120000 178.260000 13.320000 178.740000 ;
        RECT 12.120000 172.820000 13.320000 173.300000 ;
        RECT 5.560000 183.700000 7.560000 184.180000 ;
        RECT 12.120000 183.700000 13.320000 184.180000 ;
        RECT 5.560000 189.140000 7.560000 189.620000 ;
        RECT 12.120000 194.580000 13.320000 195.060000 ;
        RECT 12.120000 189.140000 13.320000 189.620000 ;
        RECT 5.560000 194.580000 7.560000 195.060000 ;
        RECT 5.560000 200.020000 7.560000 200.500000 ;
        RECT 5.560000 205.460000 7.560000 205.940000 ;
        RECT 12.120000 200.020000 13.320000 200.500000 ;
        RECT 12.120000 205.460000 13.320000 205.940000 ;
        RECT 57.120000 183.700000 58.320000 184.180000 ;
        RECT 57.120000 178.260000 58.320000 178.740000 ;
        RECT 57.120000 172.820000 58.320000 173.300000 ;
        RECT 57.120000 194.580000 58.320000 195.060000 ;
        RECT 57.120000 189.140000 58.320000 189.620000 ;
        RECT 57.120000 200.020000 58.320000 200.500000 ;
        RECT 57.120000 205.460000 58.320000 205.940000 ;
        RECT 102.120000 145.620000 103.320000 146.100000 ;
        RECT 102.120000 140.180000 103.320000 140.660000 ;
        RECT 102.120000 151.060000 103.320000 151.540000 ;
        RECT 102.120000 156.500000 103.320000 156.980000 ;
        RECT 102.120000 161.940000 103.320000 162.420000 ;
        RECT 102.120000 167.380000 103.320000 167.860000 ;
        RECT 102.120000 205.460000 103.320000 205.940000 ;
        RECT 102.120000 200.020000 103.320000 200.500000 ;
        RECT 102.120000 194.580000 103.320000 195.060000 ;
        RECT 102.120000 172.820000 103.320000 173.300000 ;
        RECT 102.120000 178.260000 103.320000 178.740000 ;
        RECT 102.120000 183.700000 103.320000 184.180000 ;
        RECT 102.120000 189.140000 103.320000 189.620000 ;
        RECT 5.560000 210.900000 7.560000 211.380000 ;
        RECT 12.120000 210.900000 13.320000 211.380000 ;
        RECT 5.560000 216.340000 7.560000 216.820000 ;
        RECT 5.560000 221.780000 7.560000 222.260000 ;
        RECT 12.120000 221.780000 13.320000 222.260000 ;
        RECT 12.120000 216.340000 13.320000 216.820000 ;
        RECT 5.560000 227.220000 7.560000 227.700000 ;
        RECT 12.120000 227.220000 13.320000 227.700000 ;
        RECT 5.560000 232.660000 7.560000 233.140000 ;
        RECT 5.560000 238.100000 7.560000 238.580000 ;
        RECT 12.120000 238.100000 13.320000 238.580000 ;
        RECT 12.120000 232.660000 13.320000 233.140000 ;
        RECT 57.120000 221.780000 58.320000 222.260000 ;
        RECT 57.120000 216.340000 58.320000 216.820000 ;
        RECT 57.120000 210.900000 58.320000 211.380000 ;
        RECT 57.120000 227.220000 58.320000 227.700000 ;
        RECT 57.120000 232.660000 58.320000 233.140000 ;
        RECT 57.120000 238.100000 58.320000 238.580000 ;
        RECT 12.120000 248.980000 13.320000 249.460000 ;
        RECT 5.560000 248.980000 7.560000 249.460000 ;
        RECT 12.120000 243.540000 13.320000 244.020000 ;
        RECT 5.560000 243.540000 7.560000 244.020000 ;
        RECT 5.560000 254.420000 7.560000 254.900000 ;
        RECT 12.120000 254.420000 13.320000 254.900000 ;
        RECT 5.560000 259.860000 7.560000 260.340000 ;
        RECT 5.560000 265.300000 7.560000 265.780000 ;
        RECT 12.120000 265.300000 13.320000 265.780000 ;
        RECT 12.120000 259.860000 13.320000 260.340000 ;
        RECT 5.560000 270.740000 7.560000 271.220000 ;
        RECT 12.120000 270.740000 13.320000 271.220000 ;
        RECT 57.120000 254.420000 58.320000 254.900000 ;
        RECT 57.120000 248.980000 58.320000 249.460000 ;
        RECT 57.120000 243.540000 58.320000 244.020000 ;
        RECT 57.120000 265.300000 58.320000 265.780000 ;
        RECT 57.120000 259.860000 58.320000 260.340000 ;
        RECT 57.120000 270.740000 58.320000 271.220000 ;
        RECT 102.120000 221.780000 103.320000 222.260000 ;
        RECT 102.120000 216.340000 103.320000 216.820000 ;
        RECT 102.120000 210.900000 103.320000 211.380000 ;
        RECT 102.120000 227.220000 103.320000 227.700000 ;
        RECT 102.120000 232.660000 103.320000 233.140000 ;
        RECT 102.120000 238.100000 103.320000 238.580000 ;
        RECT 102.120000 270.740000 103.320000 271.220000 ;
        RECT 102.120000 265.300000 103.320000 265.780000 ;
        RECT 102.120000 243.540000 103.320000 244.020000 ;
        RECT 102.120000 248.980000 103.320000 249.460000 ;
        RECT 102.120000 254.420000 103.320000 254.900000 ;
        RECT 102.120000 259.860000 103.320000 260.340000 ;
        RECT 147.120000 140.180000 148.320000 140.660000 ;
        RECT 147.120000 145.620000 148.320000 146.100000 ;
        RECT 147.120000 151.060000 148.320000 151.540000 ;
        RECT 147.120000 167.380000 148.320000 167.860000 ;
        RECT 147.120000 156.500000 148.320000 156.980000 ;
        RECT 147.120000 161.940000 148.320000 162.420000 ;
        RECT 192.120000 140.180000 193.320000 140.660000 ;
        RECT 192.120000 145.620000 193.320000 146.100000 ;
        RECT 192.120000 151.060000 193.320000 151.540000 ;
        RECT 192.120000 156.500000 193.320000 156.980000 ;
        RECT 192.120000 161.940000 193.320000 162.420000 ;
        RECT 192.120000 167.380000 193.320000 167.860000 ;
        RECT 147.120000 183.700000 148.320000 184.180000 ;
        RECT 147.120000 178.260000 148.320000 178.740000 ;
        RECT 147.120000 172.820000 148.320000 173.300000 ;
        RECT 147.120000 194.580000 148.320000 195.060000 ;
        RECT 147.120000 189.140000 148.320000 189.620000 ;
        RECT 147.120000 200.020000 148.320000 200.500000 ;
        RECT 147.120000 205.460000 148.320000 205.940000 ;
        RECT 192.120000 183.700000 193.320000 184.180000 ;
        RECT 192.120000 178.260000 193.320000 178.740000 ;
        RECT 192.120000 172.820000 193.320000 173.300000 ;
        RECT 192.120000 194.580000 193.320000 195.060000 ;
        RECT 192.120000 189.140000 193.320000 189.620000 ;
        RECT 192.120000 200.020000 193.320000 200.500000 ;
        RECT 192.120000 205.460000 193.320000 205.940000 ;
        RECT 237.120000 145.620000 238.320000 146.100000 ;
        RECT 237.120000 140.180000 238.320000 140.660000 ;
        RECT 237.120000 151.060000 238.320000 151.540000 ;
        RECT 237.120000 156.500000 238.320000 156.980000 ;
        RECT 237.120000 161.940000 238.320000 162.420000 ;
        RECT 237.120000 167.380000 238.320000 167.860000 ;
        RECT 237.120000 172.820000 238.320000 173.300000 ;
        RECT 237.120000 178.260000 238.320000 178.740000 ;
        RECT 237.120000 183.700000 238.320000 184.180000 ;
        RECT 237.120000 205.460000 238.320000 205.940000 ;
        RECT 237.120000 200.020000 238.320000 200.500000 ;
        RECT 237.120000 194.580000 238.320000 195.060000 ;
        RECT 237.120000 189.140000 238.320000 189.620000 ;
        RECT 147.120000 221.780000 148.320000 222.260000 ;
        RECT 147.120000 216.340000 148.320000 216.820000 ;
        RECT 147.120000 210.900000 148.320000 211.380000 ;
        RECT 147.120000 238.100000 148.320000 238.580000 ;
        RECT 147.120000 227.220000 148.320000 227.700000 ;
        RECT 147.120000 232.660000 148.320000 233.140000 ;
        RECT 192.120000 221.780000 193.320000 222.260000 ;
        RECT 192.120000 216.340000 193.320000 216.820000 ;
        RECT 192.120000 210.900000 193.320000 211.380000 ;
        RECT 192.120000 227.220000 193.320000 227.700000 ;
        RECT 192.120000 232.660000 193.320000 233.140000 ;
        RECT 192.120000 238.100000 193.320000 238.580000 ;
        RECT 147.120000 254.420000 148.320000 254.900000 ;
        RECT 147.120000 248.980000 148.320000 249.460000 ;
        RECT 147.120000 243.540000 148.320000 244.020000 ;
        RECT 147.120000 265.300000 148.320000 265.780000 ;
        RECT 147.120000 259.860000 148.320000 260.340000 ;
        RECT 147.120000 270.740000 148.320000 271.220000 ;
        RECT 192.120000 254.420000 193.320000 254.900000 ;
        RECT 192.120000 248.980000 193.320000 249.460000 ;
        RECT 192.120000 243.540000 193.320000 244.020000 ;
        RECT 192.120000 265.300000 193.320000 265.780000 ;
        RECT 192.120000 259.860000 193.320000 260.340000 ;
        RECT 192.120000 270.740000 193.320000 271.220000 ;
        RECT 237.120000 221.780000 238.320000 222.260000 ;
        RECT 237.120000 216.340000 238.320000 216.820000 ;
        RECT 237.120000 210.900000 238.320000 211.380000 ;
        RECT 237.120000 227.220000 238.320000 227.700000 ;
        RECT 237.120000 232.660000 238.320000 233.140000 ;
        RECT 237.120000 238.100000 238.320000 238.580000 ;
        RECT 237.120000 243.540000 238.320000 244.020000 ;
        RECT 237.120000 248.980000 238.320000 249.460000 ;
        RECT 237.120000 254.420000 238.320000 254.900000 ;
        RECT 237.120000 270.740000 238.320000 271.220000 ;
        RECT 237.120000 265.300000 238.320000 265.780000 ;
        RECT 237.120000 259.860000 238.320000 260.340000 ;
        RECT 282.120000 31.380000 283.320000 31.860000 ;
        RECT 282.120000 25.940000 283.320000 26.420000 ;
        RECT 282.120000 20.500000 283.320000 20.980000 ;
        RECT 282.120000 15.060000 283.320000 15.540000 ;
        RECT 282.120000 9.620000 283.320000 10.100000 ;
        RECT 327.120000 31.380000 328.320000 31.860000 ;
        RECT 327.120000 25.940000 328.320000 26.420000 ;
        RECT 327.120000 20.500000 328.320000 20.980000 ;
        RECT 327.120000 15.060000 328.320000 15.540000 ;
        RECT 327.120000 9.620000 328.320000 10.100000 ;
        RECT 282.120000 47.700000 283.320000 48.180000 ;
        RECT 282.120000 42.260000 283.320000 42.740000 ;
        RECT 282.120000 36.820000 283.320000 37.300000 ;
        RECT 282.120000 58.580000 283.320000 59.060000 ;
        RECT 282.120000 53.140000 283.320000 53.620000 ;
        RECT 282.120000 64.020000 283.320000 64.500000 ;
        RECT 327.120000 47.700000 328.320000 48.180000 ;
        RECT 327.120000 42.260000 328.320000 42.740000 ;
        RECT 327.120000 36.820000 328.320000 37.300000 ;
        RECT 327.120000 58.580000 328.320000 59.060000 ;
        RECT 327.120000 53.140000 328.320000 53.620000 ;
        RECT 327.120000 64.020000 328.320000 64.500000 ;
        RECT 372.120000 20.500000 373.320000 20.980000 ;
        RECT 372.120000 9.620000 373.320000 10.100000 ;
        RECT 372.120000 15.060000 373.320000 15.540000 ;
        RECT 372.120000 25.940000 373.320000 26.420000 ;
        RECT 372.120000 31.380000 373.320000 31.860000 ;
        RECT 372.120000 36.820000 373.320000 37.300000 ;
        RECT 372.120000 42.260000 373.320000 42.740000 ;
        RECT 372.120000 47.700000 373.320000 48.180000 ;
        RECT 372.120000 64.020000 373.320000 64.500000 ;
        RECT 372.120000 53.140000 373.320000 53.620000 ;
        RECT 372.120000 58.580000 373.320000 59.060000 ;
        RECT 282.120000 80.340000 283.320000 80.820000 ;
        RECT 282.120000 74.900000 283.320000 75.380000 ;
        RECT 282.120000 69.460000 283.320000 69.940000 ;
        RECT 282.120000 96.660000 283.320000 97.140000 ;
        RECT 282.120000 85.780000 283.320000 86.260000 ;
        RECT 282.120000 91.220000 283.320000 91.700000 ;
        RECT 282.120000 102.100000 283.320000 102.580000 ;
        RECT 327.120000 80.340000 328.320000 80.820000 ;
        RECT 327.120000 74.900000 328.320000 75.380000 ;
        RECT 327.120000 69.460000 328.320000 69.940000 ;
        RECT 327.120000 85.780000 328.320000 86.260000 ;
        RECT 327.120000 91.220000 328.320000 91.700000 ;
        RECT 327.120000 96.660000 328.320000 97.140000 ;
        RECT 327.120000 102.100000 328.320000 102.580000 ;
        RECT 282.120000 118.420000 283.320000 118.900000 ;
        RECT 282.120000 112.980000 283.320000 113.460000 ;
        RECT 282.120000 107.540000 283.320000 108.020000 ;
        RECT 282.120000 129.300000 283.320000 129.780000 ;
        RECT 282.120000 123.860000 283.320000 124.340000 ;
        RECT 282.120000 134.740000 283.320000 135.220000 ;
        RECT 327.120000 118.420000 328.320000 118.900000 ;
        RECT 327.120000 112.980000 328.320000 113.460000 ;
        RECT 327.120000 107.540000 328.320000 108.020000 ;
        RECT 327.120000 129.300000 328.320000 129.780000 ;
        RECT 327.120000 123.860000 328.320000 124.340000 ;
        RECT 327.120000 134.740000 328.320000 135.220000 ;
        RECT 372.120000 80.340000 373.320000 80.820000 ;
        RECT 372.120000 74.900000 373.320000 75.380000 ;
        RECT 372.120000 69.460000 373.320000 69.940000 ;
        RECT 372.120000 85.780000 373.320000 86.260000 ;
        RECT 372.120000 91.220000 373.320000 91.700000 ;
        RECT 372.120000 96.660000 373.320000 97.140000 ;
        RECT 372.120000 102.100000 373.320000 102.580000 ;
        RECT 372.120000 107.540000 373.320000 108.020000 ;
        RECT 372.120000 112.980000 373.320000 113.460000 ;
        RECT 372.120000 118.420000 373.320000 118.900000 ;
        RECT 372.120000 134.740000 373.320000 135.220000 ;
        RECT 372.120000 129.300000 373.320000 129.780000 ;
        RECT 372.120000 123.860000 373.320000 124.340000 ;
        RECT 417.120000 31.380000 418.320000 31.860000 ;
        RECT 417.120000 25.940000 418.320000 26.420000 ;
        RECT 417.120000 20.500000 418.320000 20.980000 ;
        RECT 417.120000 15.060000 418.320000 15.540000 ;
        RECT 417.120000 9.620000 418.320000 10.100000 ;
        RECT 462.120000 31.380000 463.320000 31.860000 ;
        RECT 462.120000 25.940000 463.320000 26.420000 ;
        RECT 462.120000 20.500000 463.320000 20.980000 ;
        RECT 462.120000 15.060000 463.320000 15.540000 ;
        RECT 462.120000 9.620000 463.320000 10.100000 ;
        RECT 417.120000 47.700000 418.320000 48.180000 ;
        RECT 417.120000 42.260000 418.320000 42.740000 ;
        RECT 417.120000 36.820000 418.320000 37.300000 ;
        RECT 417.120000 58.580000 418.320000 59.060000 ;
        RECT 417.120000 53.140000 418.320000 53.620000 ;
        RECT 417.120000 64.020000 418.320000 64.500000 ;
        RECT 462.120000 47.700000 463.320000 48.180000 ;
        RECT 462.120000 42.260000 463.320000 42.740000 ;
        RECT 462.120000 36.820000 463.320000 37.300000 ;
        RECT 462.120000 58.580000 463.320000 59.060000 ;
        RECT 462.120000 53.140000 463.320000 53.620000 ;
        RECT 462.120000 64.020000 463.320000 64.500000 ;
        RECT 507.120000 31.380000 508.320000 31.860000 ;
        RECT 507.120000 25.940000 508.320000 26.420000 ;
        RECT 507.120000 20.500000 508.320000 20.980000 ;
        RECT 507.120000 15.060000 508.320000 15.540000 ;
        RECT 507.120000 9.620000 508.320000 10.100000 ;
        RECT 542.600000 15.060000 544.600000 15.540000 ;
        RECT 542.600000 9.620000 544.600000 10.100000 ;
        RECT 542.600000 31.380000 544.600000 31.860000 ;
        RECT 542.600000 25.940000 544.600000 26.420000 ;
        RECT 542.600000 20.500000 544.600000 20.980000 ;
        RECT 507.120000 36.820000 508.320000 37.300000 ;
        RECT 507.120000 42.260000 508.320000 42.740000 ;
        RECT 507.120000 47.700000 508.320000 48.180000 ;
        RECT 507.120000 64.020000 508.320000 64.500000 ;
        RECT 507.120000 58.580000 508.320000 59.060000 ;
        RECT 507.120000 53.140000 508.320000 53.620000 ;
        RECT 542.600000 47.700000 544.600000 48.180000 ;
        RECT 542.600000 42.260000 544.600000 42.740000 ;
        RECT 542.600000 36.820000 544.600000 37.300000 ;
        RECT 542.600000 64.020000 544.600000 64.500000 ;
        RECT 542.600000 58.580000 544.600000 59.060000 ;
        RECT 542.600000 53.140000 544.600000 53.620000 ;
        RECT 417.120000 80.340000 418.320000 80.820000 ;
        RECT 417.120000 74.900000 418.320000 75.380000 ;
        RECT 417.120000 69.460000 418.320000 69.940000 ;
        RECT 417.120000 96.660000 418.320000 97.140000 ;
        RECT 417.120000 85.780000 418.320000 86.260000 ;
        RECT 417.120000 91.220000 418.320000 91.700000 ;
        RECT 417.120000 102.100000 418.320000 102.580000 ;
        RECT 462.120000 80.340000 463.320000 80.820000 ;
        RECT 462.120000 74.900000 463.320000 75.380000 ;
        RECT 462.120000 69.460000 463.320000 69.940000 ;
        RECT 462.120000 85.780000 463.320000 86.260000 ;
        RECT 462.120000 91.220000 463.320000 91.700000 ;
        RECT 462.120000 96.660000 463.320000 97.140000 ;
        RECT 462.120000 102.100000 463.320000 102.580000 ;
        RECT 417.120000 118.420000 418.320000 118.900000 ;
        RECT 417.120000 112.980000 418.320000 113.460000 ;
        RECT 417.120000 107.540000 418.320000 108.020000 ;
        RECT 417.120000 129.300000 418.320000 129.780000 ;
        RECT 417.120000 123.860000 418.320000 124.340000 ;
        RECT 417.120000 134.740000 418.320000 135.220000 ;
        RECT 462.120000 118.420000 463.320000 118.900000 ;
        RECT 462.120000 112.980000 463.320000 113.460000 ;
        RECT 462.120000 107.540000 463.320000 108.020000 ;
        RECT 462.120000 129.300000 463.320000 129.780000 ;
        RECT 462.120000 123.860000 463.320000 124.340000 ;
        RECT 462.120000 134.740000 463.320000 135.220000 ;
        RECT 507.120000 80.340000 508.320000 80.820000 ;
        RECT 507.120000 74.900000 508.320000 75.380000 ;
        RECT 507.120000 69.460000 508.320000 69.940000 ;
        RECT 507.120000 85.780000 508.320000 86.260000 ;
        RECT 507.120000 91.220000 508.320000 91.700000 ;
        RECT 507.120000 96.660000 508.320000 97.140000 ;
        RECT 507.120000 102.100000 508.320000 102.580000 ;
        RECT 542.600000 80.340000 544.600000 80.820000 ;
        RECT 542.600000 74.900000 544.600000 75.380000 ;
        RECT 542.600000 69.460000 544.600000 69.940000 ;
        RECT 542.600000 102.100000 544.600000 102.580000 ;
        RECT 542.600000 96.660000 544.600000 97.140000 ;
        RECT 542.600000 91.220000 544.600000 91.700000 ;
        RECT 542.600000 85.780000 544.600000 86.260000 ;
        RECT 507.120000 107.540000 508.320000 108.020000 ;
        RECT 507.120000 112.980000 508.320000 113.460000 ;
        RECT 507.120000 118.420000 508.320000 118.900000 ;
        RECT 507.120000 134.740000 508.320000 135.220000 ;
        RECT 507.120000 129.300000 508.320000 129.780000 ;
        RECT 507.120000 123.860000 508.320000 124.340000 ;
        RECT 542.600000 118.420000 544.600000 118.900000 ;
        RECT 542.600000 112.980000 544.600000 113.460000 ;
        RECT 542.600000 107.540000 544.600000 108.020000 ;
        RECT 542.600000 134.740000 544.600000 135.220000 ;
        RECT 542.600000 129.300000 544.600000 129.780000 ;
        RECT 542.600000 123.860000 544.600000 124.340000 ;
        RECT 282.120000 145.620000 283.320000 146.100000 ;
        RECT 282.120000 140.180000 283.320000 140.660000 ;
        RECT 282.120000 151.060000 283.320000 151.540000 ;
        RECT 282.120000 167.380000 283.320000 167.860000 ;
        RECT 282.120000 156.500000 283.320000 156.980000 ;
        RECT 282.120000 161.940000 283.320000 162.420000 ;
        RECT 327.120000 145.620000 328.320000 146.100000 ;
        RECT 327.120000 140.180000 328.320000 140.660000 ;
        RECT 327.120000 151.060000 328.320000 151.540000 ;
        RECT 327.120000 156.500000 328.320000 156.980000 ;
        RECT 327.120000 161.940000 328.320000 162.420000 ;
        RECT 327.120000 167.380000 328.320000 167.860000 ;
        RECT 282.120000 183.700000 283.320000 184.180000 ;
        RECT 282.120000 178.260000 283.320000 178.740000 ;
        RECT 282.120000 172.820000 283.320000 173.300000 ;
        RECT 282.120000 194.580000 283.320000 195.060000 ;
        RECT 282.120000 189.140000 283.320000 189.620000 ;
        RECT 282.120000 200.020000 283.320000 200.500000 ;
        RECT 282.120000 205.460000 283.320000 205.940000 ;
        RECT 327.120000 183.700000 328.320000 184.180000 ;
        RECT 327.120000 178.260000 328.320000 178.740000 ;
        RECT 327.120000 172.820000 328.320000 173.300000 ;
        RECT 327.120000 194.580000 328.320000 195.060000 ;
        RECT 327.120000 189.140000 328.320000 189.620000 ;
        RECT 327.120000 200.020000 328.320000 200.500000 ;
        RECT 327.120000 205.460000 328.320000 205.940000 ;
        RECT 372.120000 145.620000 373.320000 146.100000 ;
        RECT 372.120000 140.180000 373.320000 140.660000 ;
        RECT 372.120000 151.060000 373.320000 151.540000 ;
        RECT 372.120000 156.500000 373.320000 156.980000 ;
        RECT 372.120000 161.940000 373.320000 162.420000 ;
        RECT 372.120000 167.380000 373.320000 167.860000 ;
        RECT 372.120000 172.820000 373.320000 173.300000 ;
        RECT 372.120000 178.260000 373.320000 178.740000 ;
        RECT 372.120000 183.700000 373.320000 184.180000 ;
        RECT 372.120000 205.460000 373.320000 205.940000 ;
        RECT 372.120000 200.020000 373.320000 200.500000 ;
        RECT 372.120000 194.580000 373.320000 195.060000 ;
        RECT 372.120000 189.140000 373.320000 189.620000 ;
        RECT 282.120000 221.780000 283.320000 222.260000 ;
        RECT 282.120000 216.340000 283.320000 216.820000 ;
        RECT 282.120000 210.900000 283.320000 211.380000 ;
        RECT 282.120000 238.100000 283.320000 238.580000 ;
        RECT 282.120000 227.220000 283.320000 227.700000 ;
        RECT 282.120000 232.660000 283.320000 233.140000 ;
        RECT 327.120000 221.780000 328.320000 222.260000 ;
        RECT 327.120000 216.340000 328.320000 216.820000 ;
        RECT 327.120000 210.900000 328.320000 211.380000 ;
        RECT 327.120000 227.220000 328.320000 227.700000 ;
        RECT 327.120000 232.660000 328.320000 233.140000 ;
        RECT 327.120000 238.100000 328.320000 238.580000 ;
        RECT 282.120000 254.420000 283.320000 254.900000 ;
        RECT 282.120000 248.980000 283.320000 249.460000 ;
        RECT 282.120000 243.540000 283.320000 244.020000 ;
        RECT 282.120000 265.300000 283.320000 265.780000 ;
        RECT 282.120000 259.860000 283.320000 260.340000 ;
        RECT 282.120000 270.740000 283.320000 271.220000 ;
        RECT 327.120000 254.420000 328.320000 254.900000 ;
        RECT 327.120000 248.980000 328.320000 249.460000 ;
        RECT 327.120000 243.540000 328.320000 244.020000 ;
        RECT 327.120000 265.300000 328.320000 265.780000 ;
        RECT 327.120000 259.860000 328.320000 260.340000 ;
        RECT 327.120000 270.740000 328.320000 271.220000 ;
        RECT 372.120000 221.780000 373.320000 222.260000 ;
        RECT 372.120000 216.340000 373.320000 216.820000 ;
        RECT 372.120000 210.900000 373.320000 211.380000 ;
        RECT 372.120000 227.220000 373.320000 227.700000 ;
        RECT 372.120000 232.660000 373.320000 233.140000 ;
        RECT 372.120000 238.100000 373.320000 238.580000 ;
        RECT 372.120000 243.540000 373.320000 244.020000 ;
        RECT 372.120000 248.980000 373.320000 249.460000 ;
        RECT 372.120000 254.420000 373.320000 254.900000 ;
        RECT 372.120000 270.740000 373.320000 271.220000 ;
        RECT 372.120000 265.300000 373.320000 265.780000 ;
        RECT 372.120000 259.860000 373.320000 260.340000 ;
        RECT 417.120000 145.620000 418.320000 146.100000 ;
        RECT 417.120000 140.180000 418.320000 140.660000 ;
        RECT 417.120000 151.060000 418.320000 151.540000 ;
        RECT 417.120000 167.380000 418.320000 167.860000 ;
        RECT 417.120000 156.500000 418.320000 156.980000 ;
        RECT 417.120000 161.940000 418.320000 162.420000 ;
        RECT 462.120000 140.180000 463.320000 140.660000 ;
        RECT 462.120000 145.620000 463.320000 146.100000 ;
        RECT 462.120000 151.060000 463.320000 151.540000 ;
        RECT 462.120000 156.500000 463.320000 156.980000 ;
        RECT 462.120000 161.940000 463.320000 162.420000 ;
        RECT 462.120000 167.380000 463.320000 167.860000 ;
        RECT 417.120000 183.700000 418.320000 184.180000 ;
        RECT 417.120000 178.260000 418.320000 178.740000 ;
        RECT 417.120000 172.820000 418.320000 173.300000 ;
        RECT 417.120000 194.580000 418.320000 195.060000 ;
        RECT 417.120000 189.140000 418.320000 189.620000 ;
        RECT 417.120000 200.020000 418.320000 200.500000 ;
        RECT 417.120000 205.460000 418.320000 205.940000 ;
        RECT 462.120000 183.700000 463.320000 184.180000 ;
        RECT 462.120000 178.260000 463.320000 178.740000 ;
        RECT 462.120000 172.820000 463.320000 173.300000 ;
        RECT 462.120000 194.580000 463.320000 195.060000 ;
        RECT 462.120000 189.140000 463.320000 189.620000 ;
        RECT 462.120000 200.020000 463.320000 200.500000 ;
        RECT 462.120000 205.460000 463.320000 205.940000 ;
        RECT 507.120000 140.180000 508.320000 140.660000 ;
        RECT 507.120000 145.620000 508.320000 146.100000 ;
        RECT 507.120000 151.060000 508.320000 151.540000 ;
        RECT 507.120000 156.500000 508.320000 156.980000 ;
        RECT 507.120000 161.940000 508.320000 162.420000 ;
        RECT 507.120000 167.380000 508.320000 167.860000 ;
        RECT 542.600000 151.060000 544.600000 151.540000 ;
        RECT 542.600000 145.620000 544.600000 146.100000 ;
        RECT 542.600000 140.180000 544.600000 140.660000 ;
        RECT 542.600000 167.380000 544.600000 167.860000 ;
        RECT 542.600000 161.940000 544.600000 162.420000 ;
        RECT 542.600000 156.500000 544.600000 156.980000 ;
        RECT 507.120000 172.820000 508.320000 173.300000 ;
        RECT 507.120000 178.260000 508.320000 178.740000 ;
        RECT 507.120000 183.700000 508.320000 184.180000 ;
        RECT 507.120000 205.460000 508.320000 205.940000 ;
        RECT 507.120000 200.020000 508.320000 200.500000 ;
        RECT 507.120000 194.580000 508.320000 195.060000 ;
        RECT 507.120000 189.140000 508.320000 189.620000 ;
        RECT 542.600000 183.700000 544.600000 184.180000 ;
        RECT 542.600000 178.260000 544.600000 178.740000 ;
        RECT 542.600000 172.820000 544.600000 173.300000 ;
        RECT 542.600000 205.460000 544.600000 205.940000 ;
        RECT 542.600000 200.020000 544.600000 200.500000 ;
        RECT 542.600000 194.580000 544.600000 195.060000 ;
        RECT 542.600000 189.140000 544.600000 189.620000 ;
        RECT 417.120000 221.780000 418.320000 222.260000 ;
        RECT 417.120000 216.340000 418.320000 216.820000 ;
        RECT 417.120000 210.900000 418.320000 211.380000 ;
        RECT 417.120000 238.100000 418.320000 238.580000 ;
        RECT 417.120000 227.220000 418.320000 227.700000 ;
        RECT 417.120000 232.660000 418.320000 233.140000 ;
        RECT 462.120000 221.780000 463.320000 222.260000 ;
        RECT 462.120000 216.340000 463.320000 216.820000 ;
        RECT 462.120000 210.900000 463.320000 211.380000 ;
        RECT 462.120000 227.220000 463.320000 227.700000 ;
        RECT 462.120000 232.660000 463.320000 233.140000 ;
        RECT 462.120000 238.100000 463.320000 238.580000 ;
        RECT 417.120000 254.420000 418.320000 254.900000 ;
        RECT 417.120000 248.980000 418.320000 249.460000 ;
        RECT 417.120000 243.540000 418.320000 244.020000 ;
        RECT 417.120000 265.300000 418.320000 265.780000 ;
        RECT 417.120000 259.860000 418.320000 260.340000 ;
        RECT 417.120000 270.740000 418.320000 271.220000 ;
        RECT 462.120000 254.420000 463.320000 254.900000 ;
        RECT 462.120000 248.980000 463.320000 249.460000 ;
        RECT 462.120000 243.540000 463.320000 244.020000 ;
        RECT 462.120000 265.300000 463.320000 265.780000 ;
        RECT 462.120000 259.860000 463.320000 260.340000 ;
        RECT 462.120000 270.740000 463.320000 271.220000 ;
        RECT 507.120000 221.780000 508.320000 222.260000 ;
        RECT 507.120000 216.340000 508.320000 216.820000 ;
        RECT 507.120000 210.900000 508.320000 211.380000 ;
        RECT 507.120000 227.220000 508.320000 227.700000 ;
        RECT 507.120000 232.660000 508.320000 233.140000 ;
        RECT 507.120000 238.100000 508.320000 238.580000 ;
        RECT 542.600000 221.780000 544.600000 222.260000 ;
        RECT 542.600000 216.340000 544.600000 216.820000 ;
        RECT 542.600000 210.900000 544.600000 211.380000 ;
        RECT 542.600000 238.100000 544.600000 238.580000 ;
        RECT 542.600000 232.660000 544.600000 233.140000 ;
        RECT 542.600000 227.220000 544.600000 227.700000 ;
        RECT 507.120000 243.540000 508.320000 244.020000 ;
        RECT 507.120000 248.980000 508.320000 249.460000 ;
        RECT 507.120000 254.420000 508.320000 254.900000 ;
        RECT 507.120000 270.740000 508.320000 271.220000 ;
        RECT 507.120000 265.300000 508.320000 265.780000 ;
        RECT 507.120000 259.860000 508.320000 260.340000 ;
        RECT 542.600000 254.420000 544.600000 254.900000 ;
        RECT 542.600000 248.980000 544.600000 249.460000 ;
        RECT 542.600000 243.540000 544.600000 244.020000 ;
        RECT 542.600000 270.740000 544.600000 271.220000 ;
        RECT 542.600000 265.300000 544.600000 265.780000 ;
        RECT 542.600000 259.860000 544.600000 260.340000 ;
        RECT 5.560000 412.180000 7.560000 412.660000 ;
        RECT 192.120000 412.180000 193.320000 412.660000 ;
        RECT 147.120000 412.180000 148.320000 412.660000 ;
        RECT 102.120000 412.180000 103.320000 412.660000 ;
        RECT 57.120000 412.180000 58.320000 412.660000 ;
        RECT 12.120000 412.180000 13.320000 412.660000 ;
        RECT 237.120000 412.180000 238.320000 412.660000 ;
        RECT 5.560000 308.820000 7.560000 309.300000 ;
        RECT 57.120000 308.820000 58.320000 309.300000 ;
        RECT 12.120000 308.820000 13.320000 309.300000 ;
        RECT 5.560000 276.180000 7.560000 276.660000 ;
        RECT 5.560000 281.620000 7.560000 282.100000 ;
        RECT 12.120000 281.620000 13.320000 282.100000 ;
        RECT 12.120000 276.180000 13.320000 276.660000 ;
        RECT 5.560000 287.060000 7.560000 287.540000 ;
        RECT 12.120000 287.060000 13.320000 287.540000 ;
        RECT 5.560000 292.500000 7.560000 292.980000 ;
        RECT 5.560000 297.940000 7.560000 298.420000 ;
        RECT 12.120000 292.500000 13.320000 292.980000 ;
        RECT 12.120000 297.940000 13.320000 298.420000 ;
        RECT 5.560000 303.380000 7.560000 303.860000 ;
        RECT 12.120000 303.380000 13.320000 303.860000 ;
        RECT 57.120000 281.620000 58.320000 282.100000 ;
        RECT 57.120000 276.180000 58.320000 276.660000 ;
        RECT 57.120000 287.060000 58.320000 287.540000 ;
        RECT 57.120000 292.500000 58.320000 292.980000 ;
        RECT 57.120000 297.940000 58.320000 298.420000 ;
        RECT 57.120000 303.380000 58.320000 303.860000 ;
        RECT 5.560000 314.260000 7.560000 314.740000 ;
        RECT 12.120000 314.260000 13.320000 314.740000 ;
        RECT 5.560000 319.700000 7.560000 320.180000 ;
        RECT 5.560000 325.140000 7.560000 325.620000 ;
        RECT 12.120000 325.140000 13.320000 325.620000 ;
        RECT 12.120000 319.700000 13.320000 320.180000 ;
        RECT 5.560000 330.580000 7.560000 331.060000 ;
        RECT 12.120000 330.580000 13.320000 331.060000 ;
        RECT 5.560000 336.020000 7.560000 336.500000 ;
        RECT 5.560000 341.460000 7.560000 341.940000 ;
        RECT 12.120000 336.020000 13.320000 336.500000 ;
        RECT 12.120000 341.460000 13.320000 341.940000 ;
        RECT 57.120000 325.140000 58.320000 325.620000 ;
        RECT 57.120000 319.700000 58.320000 320.180000 ;
        RECT 57.120000 314.260000 58.320000 314.740000 ;
        RECT 57.120000 336.020000 58.320000 336.500000 ;
        RECT 57.120000 330.580000 58.320000 331.060000 ;
        RECT 57.120000 341.460000 58.320000 341.940000 ;
        RECT 102.120000 308.820000 103.320000 309.300000 ;
        RECT 102.120000 281.620000 103.320000 282.100000 ;
        RECT 102.120000 276.180000 103.320000 276.660000 ;
        RECT 102.120000 287.060000 103.320000 287.540000 ;
        RECT 102.120000 292.500000 103.320000 292.980000 ;
        RECT 102.120000 297.940000 103.320000 298.420000 ;
        RECT 102.120000 303.380000 103.320000 303.860000 ;
        RECT 102.120000 341.460000 103.320000 341.940000 ;
        RECT 102.120000 336.020000 103.320000 336.500000 ;
        RECT 102.120000 330.580000 103.320000 331.060000 ;
        RECT 102.120000 314.260000 103.320000 314.740000 ;
        RECT 102.120000 319.700000 103.320000 320.180000 ;
        RECT 102.120000 325.140000 103.320000 325.620000 ;
        RECT 5.560000 346.900000 7.560000 347.380000 ;
        RECT 12.120000 346.900000 13.320000 347.380000 ;
        RECT 5.560000 352.340000 7.560000 352.820000 ;
        RECT 5.560000 357.780000 7.560000 358.260000 ;
        RECT 12.120000 357.780000 13.320000 358.260000 ;
        RECT 12.120000 352.340000 13.320000 352.820000 ;
        RECT 5.560000 363.220000 7.560000 363.700000 ;
        RECT 5.560000 368.660000 7.560000 369.140000 ;
        RECT 12.120000 363.220000 13.320000 363.700000 ;
        RECT 12.120000 368.660000 13.320000 369.140000 ;
        RECT 5.560000 374.100000 7.560000 374.580000 ;
        RECT 12.120000 374.100000 13.320000 374.580000 ;
        RECT 57.120000 357.780000 58.320000 358.260000 ;
        RECT 57.120000 352.340000 58.320000 352.820000 ;
        RECT 57.120000 346.900000 58.320000 347.380000 ;
        RECT 57.120000 363.220000 58.320000 363.700000 ;
        RECT 57.120000 368.660000 58.320000 369.140000 ;
        RECT 57.120000 374.100000 58.320000 374.580000 ;
        RECT 5.560000 379.540000 7.560000 380.020000 ;
        RECT 5.560000 384.980000 7.560000 385.460000 ;
        RECT 12.120000 384.980000 13.320000 385.460000 ;
        RECT 12.120000 379.540000 13.320000 380.020000 ;
        RECT 5.560000 390.420000 7.560000 390.900000 ;
        RECT 12.120000 390.420000 13.320000 390.900000 ;
        RECT 5.560000 395.860000 7.560000 396.340000 ;
        RECT 5.560000 401.300000 7.560000 401.780000 ;
        RECT 12.120000 401.300000 13.320000 401.780000 ;
        RECT 12.120000 395.860000 13.320000 396.340000 ;
        RECT 5.560000 406.740000 7.560000 407.220000 ;
        RECT 12.120000 406.740000 13.320000 407.220000 ;
        RECT 57.120000 390.420000 58.320000 390.900000 ;
        RECT 57.120000 384.980000 58.320000 385.460000 ;
        RECT 57.120000 379.540000 58.320000 380.020000 ;
        RECT 57.120000 401.300000 58.320000 401.780000 ;
        RECT 57.120000 395.860000 58.320000 396.340000 ;
        RECT 57.120000 406.740000 58.320000 407.220000 ;
        RECT 102.120000 357.780000 103.320000 358.260000 ;
        RECT 102.120000 352.340000 103.320000 352.820000 ;
        RECT 102.120000 346.900000 103.320000 347.380000 ;
        RECT 102.120000 363.220000 103.320000 363.700000 ;
        RECT 102.120000 368.660000 103.320000 369.140000 ;
        RECT 102.120000 374.100000 103.320000 374.580000 ;
        RECT 102.120000 406.740000 103.320000 407.220000 ;
        RECT 102.120000 401.300000 103.320000 401.780000 ;
        RECT 102.120000 379.540000 103.320000 380.020000 ;
        RECT 102.120000 384.980000 103.320000 385.460000 ;
        RECT 102.120000 390.420000 103.320000 390.900000 ;
        RECT 102.120000 395.860000 103.320000 396.340000 ;
        RECT 192.120000 308.820000 193.320000 309.300000 ;
        RECT 147.120000 308.820000 148.320000 309.300000 ;
        RECT 147.120000 276.180000 148.320000 276.660000 ;
        RECT 147.120000 281.620000 148.320000 282.100000 ;
        RECT 147.120000 287.060000 148.320000 287.540000 ;
        RECT 147.120000 303.380000 148.320000 303.860000 ;
        RECT 147.120000 292.500000 148.320000 292.980000 ;
        RECT 147.120000 297.940000 148.320000 298.420000 ;
        RECT 192.120000 276.180000 193.320000 276.660000 ;
        RECT 192.120000 281.620000 193.320000 282.100000 ;
        RECT 192.120000 287.060000 193.320000 287.540000 ;
        RECT 192.120000 292.500000 193.320000 292.980000 ;
        RECT 192.120000 297.940000 193.320000 298.420000 ;
        RECT 192.120000 303.380000 193.320000 303.860000 ;
        RECT 147.120000 325.140000 148.320000 325.620000 ;
        RECT 147.120000 319.700000 148.320000 320.180000 ;
        RECT 147.120000 314.260000 148.320000 314.740000 ;
        RECT 147.120000 336.020000 148.320000 336.500000 ;
        RECT 147.120000 330.580000 148.320000 331.060000 ;
        RECT 147.120000 341.460000 148.320000 341.940000 ;
        RECT 192.120000 325.140000 193.320000 325.620000 ;
        RECT 192.120000 319.700000 193.320000 320.180000 ;
        RECT 192.120000 314.260000 193.320000 314.740000 ;
        RECT 192.120000 336.020000 193.320000 336.500000 ;
        RECT 192.120000 330.580000 193.320000 331.060000 ;
        RECT 192.120000 341.460000 193.320000 341.940000 ;
        RECT 237.120000 308.820000 238.320000 309.300000 ;
        RECT 237.120000 281.620000 238.320000 282.100000 ;
        RECT 237.120000 276.180000 238.320000 276.660000 ;
        RECT 237.120000 287.060000 238.320000 287.540000 ;
        RECT 237.120000 292.500000 238.320000 292.980000 ;
        RECT 237.120000 297.940000 238.320000 298.420000 ;
        RECT 237.120000 303.380000 238.320000 303.860000 ;
        RECT 237.120000 314.260000 238.320000 314.740000 ;
        RECT 237.120000 319.700000 238.320000 320.180000 ;
        RECT 237.120000 325.140000 238.320000 325.620000 ;
        RECT 237.120000 341.460000 238.320000 341.940000 ;
        RECT 237.120000 336.020000 238.320000 336.500000 ;
        RECT 237.120000 330.580000 238.320000 331.060000 ;
        RECT 147.120000 357.780000 148.320000 358.260000 ;
        RECT 147.120000 352.340000 148.320000 352.820000 ;
        RECT 147.120000 346.900000 148.320000 347.380000 ;
        RECT 147.120000 374.100000 148.320000 374.580000 ;
        RECT 147.120000 363.220000 148.320000 363.700000 ;
        RECT 147.120000 368.660000 148.320000 369.140000 ;
        RECT 192.120000 357.780000 193.320000 358.260000 ;
        RECT 192.120000 352.340000 193.320000 352.820000 ;
        RECT 192.120000 346.900000 193.320000 347.380000 ;
        RECT 192.120000 363.220000 193.320000 363.700000 ;
        RECT 192.120000 368.660000 193.320000 369.140000 ;
        RECT 192.120000 374.100000 193.320000 374.580000 ;
        RECT 147.120000 390.420000 148.320000 390.900000 ;
        RECT 147.120000 384.980000 148.320000 385.460000 ;
        RECT 147.120000 379.540000 148.320000 380.020000 ;
        RECT 147.120000 401.300000 148.320000 401.780000 ;
        RECT 147.120000 395.860000 148.320000 396.340000 ;
        RECT 147.120000 406.740000 148.320000 407.220000 ;
        RECT 192.120000 390.420000 193.320000 390.900000 ;
        RECT 192.120000 384.980000 193.320000 385.460000 ;
        RECT 192.120000 379.540000 193.320000 380.020000 ;
        RECT 192.120000 401.300000 193.320000 401.780000 ;
        RECT 192.120000 395.860000 193.320000 396.340000 ;
        RECT 192.120000 406.740000 193.320000 407.220000 ;
        RECT 237.120000 357.780000 238.320000 358.260000 ;
        RECT 237.120000 352.340000 238.320000 352.820000 ;
        RECT 237.120000 346.900000 238.320000 347.380000 ;
        RECT 237.120000 363.220000 238.320000 363.700000 ;
        RECT 237.120000 368.660000 238.320000 369.140000 ;
        RECT 237.120000 374.100000 238.320000 374.580000 ;
        RECT 237.120000 379.540000 238.320000 380.020000 ;
        RECT 237.120000 384.980000 238.320000 385.460000 ;
        RECT 237.120000 390.420000 238.320000 390.900000 ;
        RECT 237.120000 406.740000 238.320000 407.220000 ;
        RECT 237.120000 401.300000 238.320000 401.780000 ;
        RECT 237.120000 395.860000 238.320000 396.340000 ;
        RECT 5.560000 417.620000 7.560000 418.100000 ;
        RECT 12.120000 417.620000 13.320000 418.100000 ;
        RECT 5.560000 423.060000 7.560000 423.540000 ;
        RECT 5.560000 428.500000 7.560000 428.980000 ;
        RECT 12.120000 423.060000 13.320000 423.540000 ;
        RECT 12.120000 428.500000 13.320000 428.980000 ;
        RECT 5.560000 433.940000 7.560000 434.420000 ;
        RECT 12.120000 433.940000 13.320000 434.420000 ;
        RECT 5.560000 439.380000 7.560000 439.860000 ;
        RECT 5.560000 444.820000 7.560000 445.300000 ;
        RECT 12.120000 444.820000 13.320000 445.300000 ;
        RECT 12.120000 439.380000 13.320000 439.860000 ;
        RECT 57.120000 417.620000 58.320000 418.100000 ;
        RECT 57.120000 423.060000 58.320000 423.540000 ;
        RECT 57.120000 428.500000 58.320000 428.980000 ;
        RECT 57.120000 433.940000 58.320000 434.420000 ;
        RECT 57.120000 439.380000 58.320000 439.860000 ;
        RECT 57.120000 444.820000 58.320000 445.300000 ;
        RECT 5.560000 450.260000 7.560000 450.740000 ;
        RECT 12.120000 450.260000 13.320000 450.740000 ;
        RECT 5.560000 455.700000 7.560000 456.180000 ;
        RECT 5.560000 461.140000 7.560000 461.620000 ;
        RECT 12.120000 461.140000 13.320000 461.620000 ;
        RECT 12.120000 455.700000 13.320000 456.180000 ;
        RECT 5.560000 466.580000 7.560000 467.060000 ;
        RECT 5.560000 472.020000 7.560000 472.500000 ;
        RECT 12.120000 472.020000 13.320000 472.500000 ;
        RECT 12.120000 466.580000 13.320000 467.060000 ;
        RECT 5.560000 477.460000 7.560000 477.940000 ;
        RECT 12.120000 477.460000 13.320000 477.940000 ;
        RECT 57.120000 461.140000 58.320000 461.620000 ;
        RECT 57.120000 455.700000 58.320000 456.180000 ;
        RECT 57.120000 450.260000 58.320000 450.740000 ;
        RECT 57.120000 472.020000 58.320000 472.500000 ;
        RECT 57.120000 466.580000 58.320000 467.060000 ;
        RECT 57.120000 477.460000 58.320000 477.940000 ;
        RECT 102.120000 428.500000 103.320000 428.980000 ;
        RECT 102.120000 417.620000 103.320000 418.100000 ;
        RECT 102.120000 423.060000 103.320000 423.540000 ;
        RECT 102.120000 433.940000 103.320000 434.420000 ;
        RECT 102.120000 439.380000 103.320000 439.860000 ;
        RECT 102.120000 444.820000 103.320000 445.300000 ;
        RECT 102.120000 477.460000 103.320000 477.940000 ;
        RECT 102.120000 472.020000 103.320000 472.500000 ;
        RECT 102.120000 450.260000 103.320000 450.740000 ;
        RECT 102.120000 455.700000 103.320000 456.180000 ;
        RECT 102.120000 461.140000 103.320000 461.620000 ;
        RECT 102.120000 466.580000 103.320000 467.060000 ;
        RECT 5.560000 515.540000 7.560000 516.020000 ;
        RECT 57.120000 515.540000 58.320000 516.020000 ;
        RECT 12.120000 515.540000 13.320000 516.020000 ;
        RECT 5.560000 482.900000 7.560000 483.380000 ;
        RECT 5.560000 488.340000 7.560000 488.820000 ;
        RECT 12.120000 488.340000 13.320000 488.820000 ;
        RECT 12.120000 482.900000 13.320000 483.380000 ;
        RECT 5.560000 493.780000 7.560000 494.260000 ;
        RECT 12.120000 493.780000 13.320000 494.260000 ;
        RECT 5.560000 499.220000 7.560000 499.700000 ;
        RECT 5.560000 504.660000 7.560000 505.140000 ;
        RECT 12.120000 504.660000 13.320000 505.140000 ;
        RECT 12.120000 499.220000 13.320000 499.700000 ;
        RECT 5.560000 510.100000 7.560000 510.580000 ;
        RECT 12.120000 510.100000 13.320000 510.580000 ;
        RECT 57.120000 493.780000 58.320000 494.260000 ;
        RECT 57.120000 488.340000 58.320000 488.820000 ;
        RECT 57.120000 482.900000 58.320000 483.380000 ;
        RECT 57.120000 504.660000 58.320000 505.140000 ;
        RECT 57.120000 499.220000 58.320000 499.700000 ;
        RECT 57.120000 510.100000 58.320000 510.580000 ;
        RECT 5.560000 520.980000 7.560000 521.460000 ;
        RECT 12.120000 520.980000 13.320000 521.460000 ;
        RECT 5.560000 526.420000 7.560000 526.900000 ;
        RECT 5.560000 531.860000 7.560000 532.340000 ;
        RECT 12.120000 531.860000 13.320000 532.340000 ;
        RECT 12.120000 526.420000 13.320000 526.900000 ;
        RECT 12.120000 537.300000 13.320000 537.780000 ;
        RECT 5.560000 537.300000 7.560000 537.780000 ;
        RECT 57.120000 520.980000 58.320000 521.460000 ;
        RECT 57.120000 526.420000 58.320000 526.900000 ;
        RECT 57.120000 531.860000 58.320000 532.340000 ;
        RECT 57.120000 537.300000 58.320000 537.780000 ;
        RECT 102.120000 515.540000 103.320000 516.020000 ;
        RECT 102.120000 488.340000 103.320000 488.820000 ;
        RECT 102.120000 482.900000 103.320000 483.380000 ;
        RECT 102.120000 493.780000 103.320000 494.260000 ;
        RECT 102.120000 499.220000 103.320000 499.700000 ;
        RECT 102.120000 504.660000 103.320000 505.140000 ;
        RECT 102.120000 510.100000 103.320000 510.580000 ;
        RECT 102.120000 537.300000 103.320000 537.780000 ;
        RECT 102.120000 520.980000 103.320000 521.460000 ;
        RECT 102.120000 526.420000 103.320000 526.900000 ;
        RECT 102.120000 531.860000 103.320000 532.340000 ;
        RECT 147.120000 417.620000 148.320000 418.100000 ;
        RECT 147.120000 423.060000 148.320000 423.540000 ;
        RECT 147.120000 428.500000 148.320000 428.980000 ;
        RECT 147.120000 444.820000 148.320000 445.300000 ;
        RECT 147.120000 433.940000 148.320000 434.420000 ;
        RECT 147.120000 439.380000 148.320000 439.860000 ;
        RECT 192.120000 428.500000 193.320000 428.980000 ;
        RECT 192.120000 417.620000 193.320000 418.100000 ;
        RECT 192.120000 423.060000 193.320000 423.540000 ;
        RECT 192.120000 433.940000 193.320000 434.420000 ;
        RECT 192.120000 439.380000 193.320000 439.860000 ;
        RECT 192.120000 444.820000 193.320000 445.300000 ;
        RECT 147.120000 461.140000 148.320000 461.620000 ;
        RECT 147.120000 455.700000 148.320000 456.180000 ;
        RECT 147.120000 450.260000 148.320000 450.740000 ;
        RECT 147.120000 472.020000 148.320000 472.500000 ;
        RECT 147.120000 466.580000 148.320000 467.060000 ;
        RECT 147.120000 477.460000 148.320000 477.940000 ;
        RECT 192.120000 461.140000 193.320000 461.620000 ;
        RECT 192.120000 455.700000 193.320000 456.180000 ;
        RECT 192.120000 450.260000 193.320000 450.740000 ;
        RECT 192.120000 472.020000 193.320000 472.500000 ;
        RECT 192.120000 466.580000 193.320000 467.060000 ;
        RECT 192.120000 477.460000 193.320000 477.940000 ;
        RECT 237.120000 417.620000 238.320000 418.100000 ;
        RECT 237.120000 423.060000 238.320000 423.540000 ;
        RECT 237.120000 428.500000 238.320000 428.980000 ;
        RECT 237.120000 433.940000 238.320000 434.420000 ;
        RECT 237.120000 439.380000 238.320000 439.860000 ;
        RECT 237.120000 444.820000 238.320000 445.300000 ;
        RECT 237.120000 450.260000 238.320000 450.740000 ;
        RECT 237.120000 455.700000 238.320000 456.180000 ;
        RECT 237.120000 461.140000 238.320000 461.620000 ;
        RECT 237.120000 477.460000 238.320000 477.940000 ;
        RECT 237.120000 472.020000 238.320000 472.500000 ;
        RECT 237.120000 466.580000 238.320000 467.060000 ;
        RECT 192.120000 515.540000 193.320000 516.020000 ;
        RECT 147.120000 515.540000 148.320000 516.020000 ;
        RECT 147.120000 493.780000 148.320000 494.260000 ;
        RECT 147.120000 488.340000 148.320000 488.820000 ;
        RECT 147.120000 482.900000 148.320000 483.380000 ;
        RECT 147.120000 499.220000 148.320000 499.700000 ;
        RECT 147.120000 504.660000 148.320000 505.140000 ;
        RECT 147.120000 510.100000 148.320000 510.580000 ;
        RECT 192.120000 488.340000 193.320000 488.820000 ;
        RECT 192.120000 482.900000 193.320000 483.380000 ;
        RECT 192.120000 493.780000 193.320000 494.260000 ;
        RECT 192.120000 504.660000 193.320000 505.140000 ;
        RECT 192.120000 499.220000 193.320000 499.700000 ;
        RECT 192.120000 510.100000 193.320000 510.580000 ;
        RECT 147.120000 520.980000 148.320000 521.460000 ;
        RECT 147.120000 526.420000 148.320000 526.900000 ;
        RECT 147.120000 531.860000 148.320000 532.340000 ;
        RECT 147.120000 537.300000 148.320000 537.780000 ;
        RECT 192.120000 520.980000 193.320000 521.460000 ;
        RECT 192.120000 526.420000 193.320000 526.900000 ;
        RECT 192.120000 531.860000 193.320000 532.340000 ;
        RECT 192.120000 537.300000 193.320000 537.780000 ;
        RECT 237.120000 515.540000 238.320000 516.020000 ;
        RECT 237.120000 493.780000 238.320000 494.260000 ;
        RECT 237.120000 488.340000 238.320000 488.820000 ;
        RECT 237.120000 482.900000 238.320000 483.380000 ;
        RECT 237.120000 499.220000 238.320000 499.700000 ;
        RECT 237.120000 504.660000 238.320000 505.140000 ;
        RECT 237.120000 510.100000 238.320000 510.580000 ;
        RECT 237.120000 537.300000 238.320000 537.780000 ;
        RECT 237.120000 520.980000 238.320000 521.460000 ;
        RECT 237.120000 526.420000 238.320000 526.900000 ;
        RECT 237.120000 531.860000 238.320000 532.340000 ;
        RECT 542.600000 412.180000 544.600000 412.660000 ;
        RECT 507.120000 412.180000 508.320000 412.660000 ;
        RECT 462.120000 412.180000 463.320000 412.660000 ;
        RECT 417.120000 412.180000 418.320000 412.660000 ;
        RECT 372.120000 412.180000 373.320000 412.660000 ;
        RECT 327.120000 412.180000 328.320000 412.660000 ;
        RECT 282.120000 412.180000 283.320000 412.660000 ;
        RECT 327.120000 308.820000 328.320000 309.300000 ;
        RECT 282.120000 308.820000 283.320000 309.300000 ;
        RECT 282.120000 281.620000 283.320000 282.100000 ;
        RECT 282.120000 276.180000 283.320000 276.660000 ;
        RECT 282.120000 287.060000 283.320000 287.540000 ;
        RECT 282.120000 303.380000 283.320000 303.860000 ;
        RECT 282.120000 292.500000 283.320000 292.980000 ;
        RECT 282.120000 297.940000 283.320000 298.420000 ;
        RECT 327.120000 281.620000 328.320000 282.100000 ;
        RECT 327.120000 276.180000 328.320000 276.660000 ;
        RECT 327.120000 287.060000 328.320000 287.540000 ;
        RECT 327.120000 292.500000 328.320000 292.980000 ;
        RECT 327.120000 297.940000 328.320000 298.420000 ;
        RECT 327.120000 303.380000 328.320000 303.860000 ;
        RECT 282.120000 325.140000 283.320000 325.620000 ;
        RECT 282.120000 319.700000 283.320000 320.180000 ;
        RECT 282.120000 314.260000 283.320000 314.740000 ;
        RECT 282.120000 336.020000 283.320000 336.500000 ;
        RECT 282.120000 330.580000 283.320000 331.060000 ;
        RECT 282.120000 341.460000 283.320000 341.940000 ;
        RECT 327.120000 325.140000 328.320000 325.620000 ;
        RECT 327.120000 319.700000 328.320000 320.180000 ;
        RECT 327.120000 314.260000 328.320000 314.740000 ;
        RECT 327.120000 336.020000 328.320000 336.500000 ;
        RECT 327.120000 330.580000 328.320000 331.060000 ;
        RECT 327.120000 341.460000 328.320000 341.940000 ;
        RECT 372.120000 308.820000 373.320000 309.300000 ;
        RECT 372.120000 281.620000 373.320000 282.100000 ;
        RECT 372.120000 276.180000 373.320000 276.660000 ;
        RECT 372.120000 287.060000 373.320000 287.540000 ;
        RECT 372.120000 292.500000 373.320000 292.980000 ;
        RECT 372.120000 297.940000 373.320000 298.420000 ;
        RECT 372.120000 303.380000 373.320000 303.860000 ;
        RECT 372.120000 314.260000 373.320000 314.740000 ;
        RECT 372.120000 319.700000 373.320000 320.180000 ;
        RECT 372.120000 325.140000 373.320000 325.620000 ;
        RECT 372.120000 341.460000 373.320000 341.940000 ;
        RECT 372.120000 336.020000 373.320000 336.500000 ;
        RECT 372.120000 330.580000 373.320000 331.060000 ;
        RECT 282.120000 357.780000 283.320000 358.260000 ;
        RECT 282.120000 352.340000 283.320000 352.820000 ;
        RECT 282.120000 346.900000 283.320000 347.380000 ;
        RECT 282.120000 374.100000 283.320000 374.580000 ;
        RECT 282.120000 363.220000 283.320000 363.700000 ;
        RECT 282.120000 368.660000 283.320000 369.140000 ;
        RECT 327.120000 357.780000 328.320000 358.260000 ;
        RECT 327.120000 352.340000 328.320000 352.820000 ;
        RECT 327.120000 346.900000 328.320000 347.380000 ;
        RECT 327.120000 363.220000 328.320000 363.700000 ;
        RECT 327.120000 368.660000 328.320000 369.140000 ;
        RECT 327.120000 374.100000 328.320000 374.580000 ;
        RECT 282.120000 390.420000 283.320000 390.900000 ;
        RECT 282.120000 384.980000 283.320000 385.460000 ;
        RECT 282.120000 379.540000 283.320000 380.020000 ;
        RECT 282.120000 401.300000 283.320000 401.780000 ;
        RECT 282.120000 395.860000 283.320000 396.340000 ;
        RECT 282.120000 406.740000 283.320000 407.220000 ;
        RECT 327.120000 390.420000 328.320000 390.900000 ;
        RECT 327.120000 384.980000 328.320000 385.460000 ;
        RECT 327.120000 379.540000 328.320000 380.020000 ;
        RECT 327.120000 401.300000 328.320000 401.780000 ;
        RECT 327.120000 395.860000 328.320000 396.340000 ;
        RECT 327.120000 406.740000 328.320000 407.220000 ;
        RECT 372.120000 357.780000 373.320000 358.260000 ;
        RECT 372.120000 352.340000 373.320000 352.820000 ;
        RECT 372.120000 346.900000 373.320000 347.380000 ;
        RECT 372.120000 363.220000 373.320000 363.700000 ;
        RECT 372.120000 368.660000 373.320000 369.140000 ;
        RECT 372.120000 374.100000 373.320000 374.580000 ;
        RECT 372.120000 379.540000 373.320000 380.020000 ;
        RECT 372.120000 384.980000 373.320000 385.460000 ;
        RECT 372.120000 390.420000 373.320000 390.900000 ;
        RECT 372.120000 406.740000 373.320000 407.220000 ;
        RECT 372.120000 401.300000 373.320000 401.780000 ;
        RECT 372.120000 395.860000 373.320000 396.340000 ;
        RECT 462.120000 308.820000 463.320000 309.300000 ;
        RECT 417.120000 308.820000 418.320000 309.300000 ;
        RECT 417.120000 281.620000 418.320000 282.100000 ;
        RECT 417.120000 276.180000 418.320000 276.660000 ;
        RECT 417.120000 287.060000 418.320000 287.540000 ;
        RECT 417.120000 303.380000 418.320000 303.860000 ;
        RECT 417.120000 292.500000 418.320000 292.980000 ;
        RECT 417.120000 297.940000 418.320000 298.420000 ;
        RECT 462.120000 276.180000 463.320000 276.660000 ;
        RECT 462.120000 281.620000 463.320000 282.100000 ;
        RECT 462.120000 287.060000 463.320000 287.540000 ;
        RECT 462.120000 292.500000 463.320000 292.980000 ;
        RECT 462.120000 297.940000 463.320000 298.420000 ;
        RECT 462.120000 303.380000 463.320000 303.860000 ;
        RECT 417.120000 325.140000 418.320000 325.620000 ;
        RECT 417.120000 319.700000 418.320000 320.180000 ;
        RECT 417.120000 314.260000 418.320000 314.740000 ;
        RECT 417.120000 336.020000 418.320000 336.500000 ;
        RECT 417.120000 330.580000 418.320000 331.060000 ;
        RECT 417.120000 341.460000 418.320000 341.940000 ;
        RECT 462.120000 325.140000 463.320000 325.620000 ;
        RECT 462.120000 319.700000 463.320000 320.180000 ;
        RECT 462.120000 314.260000 463.320000 314.740000 ;
        RECT 462.120000 336.020000 463.320000 336.500000 ;
        RECT 462.120000 330.580000 463.320000 331.060000 ;
        RECT 462.120000 341.460000 463.320000 341.940000 ;
        RECT 542.600000 308.820000 544.600000 309.300000 ;
        RECT 507.120000 308.820000 508.320000 309.300000 ;
        RECT 507.120000 276.180000 508.320000 276.660000 ;
        RECT 507.120000 281.620000 508.320000 282.100000 ;
        RECT 507.120000 287.060000 508.320000 287.540000 ;
        RECT 507.120000 292.500000 508.320000 292.980000 ;
        RECT 507.120000 297.940000 508.320000 298.420000 ;
        RECT 507.120000 303.380000 508.320000 303.860000 ;
        RECT 542.600000 287.060000 544.600000 287.540000 ;
        RECT 542.600000 281.620000 544.600000 282.100000 ;
        RECT 542.600000 276.180000 544.600000 276.660000 ;
        RECT 542.600000 303.380000 544.600000 303.860000 ;
        RECT 542.600000 297.940000 544.600000 298.420000 ;
        RECT 542.600000 292.500000 544.600000 292.980000 ;
        RECT 507.120000 314.260000 508.320000 314.740000 ;
        RECT 507.120000 319.700000 508.320000 320.180000 ;
        RECT 507.120000 325.140000 508.320000 325.620000 ;
        RECT 507.120000 341.460000 508.320000 341.940000 ;
        RECT 507.120000 336.020000 508.320000 336.500000 ;
        RECT 507.120000 330.580000 508.320000 331.060000 ;
        RECT 542.600000 325.140000 544.600000 325.620000 ;
        RECT 542.600000 319.700000 544.600000 320.180000 ;
        RECT 542.600000 314.260000 544.600000 314.740000 ;
        RECT 542.600000 341.460000 544.600000 341.940000 ;
        RECT 542.600000 336.020000 544.600000 336.500000 ;
        RECT 542.600000 330.580000 544.600000 331.060000 ;
        RECT 417.120000 357.780000 418.320000 358.260000 ;
        RECT 417.120000 352.340000 418.320000 352.820000 ;
        RECT 417.120000 346.900000 418.320000 347.380000 ;
        RECT 417.120000 374.100000 418.320000 374.580000 ;
        RECT 417.120000 363.220000 418.320000 363.700000 ;
        RECT 417.120000 368.660000 418.320000 369.140000 ;
        RECT 462.120000 357.780000 463.320000 358.260000 ;
        RECT 462.120000 352.340000 463.320000 352.820000 ;
        RECT 462.120000 346.900000 463.320000 347.380000 ;
        RECT 462.120000 363.220000 463.320000 363.700000 ;
        RECT 462.120000 368.660000 463.320000 369.140000 ;
        RECT 462.120000 374.100000 463.320000 374.580000 ;
        RECT 417.120000 390.420000 418.320000 390.900000 ;
        RECT 417.120000 384.980000 418.320000 385.460000 ;
        RECT 417.120000 379.540000 418.320000 380.020000 ;
        RECT 417.120000 401.300000 418.320000 401.780000 ;
        RECT 417.120000 395.860000 418.320000 396.340000 ;
        RECT 417.120000 406.740000 418.320000 407.220000 ;
        RECT 462.120000 390.420000 463.320000 390.900000 ;
        RECT 462.120000 384.980000 463.320000 385.460000 ;
        RECT 462.120000 379.540000 463.320000 380.020000 ;
        RECT 462.120000 401.300000 463.320000 401.780000 ;
        RECT 462.120000 395.860000 463.320000 396.340000 ;
        RECT 462.120000 406.740000 463.320000 407.220000 ;
        RECT 507.120000 357.780000 508.320000 358.260000 ;
        RECT 507.120000 352.340000 508.320000 352.820000 ;
        RECT 507.120000 346.900000 508.320000 347.380000 ;
        RECT 507.120000 363.220000 508.320000 363.700000 ;
        RECT 507.120000 368.660000 508.320000 369.140000 ;
        RECT 507.120000 374.100000 508.320000 374.580000 ;
        RECT 542.600000 357.780000 544.600000 358.260000 ;
        RECT 542.600000 352.340000 544.600000 352.820000 ;
        RECT 542.600000 346.900000 544.600000 347.380000 ;
        RECT 542.600000 374.100000 544.600000 374.580000 ;
        RECT 542.600000 368.660000 544.600000 369.140000 ;
        RECT 542.600000 363.220000 544.600000 363.700000 ;
        RECT 507.120000 379.540000 508.320000 380.020000 ;
        RECT 507.120000 384.980000 508.320000 385.460000 ;
        RECT 507.120000 390.420000 508.320000 390.900000 ;
        RECT 507.120000 406.740000 508.320000 407.220000 ;
        RECT 507.120000 401.300000 508.320000 401.780000 ;
        RECT 507.120000 395.860000 508.320000 396.340000 ;
        RECT 542.600000 390.420000 544.600000 390.900000 ;
        RECT 542.600000 384.980000 544.600000 385.460000 ;
        RECT 542.600000 379.540000 544.600000 380.020000 ;
        RECT 542.600000 406.740000 544.600000 407.220000 ;
        RECT 542.600000 401.300000 544.600000 401.780000 ;
        RECT 542.600000 395.860000 544.600000 396.340000 ;
        RECT 282.120000 417.620000 283.320000 418.100000 ;
        RECT 282.120000 423.060000 283.320000 423.540000 ;
        RECT 282.120000 428.500000 283.320000 428.980000 ;
        RECT 282.120000 444.820000 283.320000 445.300000 ;
        RECT 282.120000 433.940000 283.320000 434.420000 ;
        RECT 282.120000 439.380000 283.320000 439.860000 ;
        RECT 327.120000 417.620000 328.320000 418.100000 ;
        RECT 327.120000 423.060000 328.320000 423.540000 ;
        RECT 327.120000 428.500000 328.320000 428.980000 ;
        RECT 327.120000 433.940000 328.320000 434.420000 ;
        RECT 327.120000 439.380000 328.320000 439.860000 ;
        RECT 327.120000 444.820000 328.320000 445.300000 ;
        RECT 282.120000 461.140000 283.320000 461.620000 ;
        RECT 282.120000 455.700000 283.320000 456.180000 ;
        RECT 282.120000 450.260000 283.320000 450.740000 ;
        RECT 282.120000 472.020000 283.320000 472.500000 ;
        RECT 282.120000 466.580000 283.320000 467.060000 ;
        RECT 282.120000 477.460000 283.320000 477.940000 ;
        RECT 327.120000 461.140000 328.320000 461.620000 ;
        RECT 327.120000 455.700000 328.320000 456.180000 ;
        RECT 327.120000 450.260000 328.320000 450.740000 ;
        RECT 327.120000 472.020000 328.320000 472.500000 ;
        RECT 327.120000 466.580000 328.320000 467.060000 ;
        RECT 327.120000 477.460000 328.320000 477.940000 ;
        RECT 372.120000 428.500000 373.320000 428.980000 ;
        RECT 372.120000 417.620000 373.320000 418.100000 ;
        RECT 372.120000 423.060000 373.320000 423.540000 ;
        RECT 372.120000 433.940000 373.320000 434.420000 ;
        RECT 372.120000 439.380000 373.320000 439.860000 ;
        RECT 372.120000 444.820000 373.320000 445.300000 ;
        RECT 372.120000 450.260000 373.320000 450.740000 ;
        RECT 372.120000 455.700000 373.320000 456.180000 ;
        RECT 372.120000 461.140000 373.320000 461.620000 ;
        RECT 372.120000 477.460000 373.320000 477.940000 ;
        RECT 372.120000 472.020000 373.320000 472.500000 ;
        RECT 372.120000 466.580000 373.320000 467.060000 ;
        RECT 327.120000 515.540000 328.320000 516.020000 ;
        RECT 282.120000 515.540000 283.320000 516.020000 ;
        RECT 282.120000 493.780000 283.320000 494.260000 ;
        RECT 282.120000 488.340000 283.320000 488.820000 ;
        RECT 282.120000 482.900000 283.320000 483.380000 ;
        RECT 282.120000 499.220000 283.320000 499.700000 ;
        RECT 282.120000 504.660000 283.320000 505.140000 ;
        RECT 282.120000 510.100000 283.320000 510.580000 ;
        RECT 327.120000 493.780000 328.320000 494.260000 ;
        RECT 327.120000 488.340000 328.320000 488.820000 ;
        RECT 327.120000 482.900000 328.320000 483.380000 ;
        RECT 327.120000 504.660000 328.320000 505.140000 ;
        RECT 327.120000 499.220000 328.320000 499.700000 ;
        RECT 327.120000 510.100000 328.320000 510.580000 ;
        RECT 282.120000 520.980000 283.320000 521.460000 ;
        RECT 282.120000 526.420000 283.320000 526.900000 ;
        RECT 282.120000 531.860000 283.320000 532.340000 ;
        RECT 282.120000 537.300000 283.320000 537.780000 ;
        RECT 327.120000 520.980000 328.320000 521.460000 ;
        RECT 327.120000 526.420000 328.320000 526.900000 ;
        RECT 327.120000 531.860000 328.320000 532.340000 ;
        RECT 327.120000 537.300000 328.320000 537.780000 ;
        RECT 372.120000 515.540000 373.320000 516.020000 ;
        RECT 372.120000 488.340000 373.320000 488.820000 ;
        RECT 372.120000 482.900000 373.320000 483.380000 ;
        RECT 372.120000 493.780000 373.320000 494.260000 ;
        RECT 372.120000 499.220000 373.320000 499.700000 ;
        RECT 372.120000 504.660000 373.320000 505.140000 ;
        RECT 372.120000 510.100000 373.320000 510.580000 ;
        RECT 372.120000 537.300000 373.320000 537.780000 ;
        RECT 372.120000 520.980000 373.320000 521.460000 ;
        RECT 372.120000 526.420000 373.320000 526.900000 ;
        RECT 372.120000 531.860000 373.320000 532.340000 ;
        RECT 417.120000 417.620000 418.320000 418.100000 ;
        RECT 417.120000 423.060000 418.320000 423.540000 ;
        RECT 417.120000 428.500000 418.320000 428.980000 ;
        RECT 417.120000 444.820000 418.320000 445.300000 ;
        RECT 417.120000 433.940000 418.320000 434.420000 ;
        RECT 417.120000 439.380000 418.320000 439.860000 ;
        RECT 462.120000 417.620000 463.320000 418.100000 ;
        RECT 462.120000 423.060000 463.320000 423.540000 ;
        RECT 462.120000 428.500000 463.320000 428.980000 ;
        RECT 462.120000 433.940000 463.320000 434.420000 ;
        RECT 462.120000 439.380000 463.320000 439.860000 ;
        RECT 462.120000 444.820000 463.320000 445.300000 ;
        RECT 417.120000 461.140000 418.320000 461.620000 ;
        RECT 417.120000 455.700000 418.320000 456.180000 ;
        RECT 417.120000 450.260000 418.320000 450.740000 ;
        RECT 417.120000 472.020000 418.320000 472.500000 ;
        RECT 417.120000 466.580000 418.320000 467.060000 ;
        RECT 417.120000 477.460000 418.320000 477.940000 ;
        RECT 462.120000 461.140000 463.320000 461.620000 ;
        RECT 462.120000 455.700000 463.320000 456.180000 ;
        RECT 462.120000 450.260000 463.320000 450.740000 ;
        RECT 462.120000 472.020000 463.320000 472.500000 ;
        RECT 462.120000 466.580000 463.320000 467.060000 ;
        RECT 462.120000 477.460000 463.320000 477.940000 ;
        RECT 507.120000 428.500000 508.320000 428.980000 ;
        RECT 507.120000 417.620000 508.320000 418.100000 ;
        RECT 507.120000 423.060000 508.320000 423.540000 ;
        RECT 507.120000 433.940000 508.320000 434.420000 ;
        RECT 507.120000 439.380000 508.320000 439.860000 ;
        RECT 507.120000 444.820000 508.320000 445.300000 ;
        RECT 542.600000 428.500000 544.600000 428.980000 ;
        RECT 542.600000 423.060000 544.600000 423.540000 ;
        RECT 542.600000 417.620000 544.600000 418.100000 ;
        RECT 542.600000 444.820000 544.600000 445.300000 ;
        RECT 542.600000 439.380000 544.600000 439.860000 ;
        RECT 542.600000 433.940000 544.600000 434.420000 ;
        RECT 507.120000 450.260000 508.320000 450.740000 ;
        RECT 507.120000 455.700000 508.320000 456.180000 ;
        RECT 507.120000 461.140000 508.320000 461.620000 ;
        RECT 507.120000 477.460000 508.320000 477.940000 ;
        RECT 507.120000 472.020000 508.320000 472.500000 ;
        RECT 507.120000 466.580000 508.320000 467.060000 ;
        RECT 542.600000 461.140000 544.600000 461.620000 ;
        RECT 542.600000 455.700000 544.600000 456.180000 ;
        RECT 542.600000 450.260000 544.600000 450.740000 ;
        RECT 542.600000 477.460000 544.600000 477.940000 ;
        RECT 542.600000 472.020000 544.600000 472.500000 ;
        RECT 542.600000 466.580000 544.600000 467.060000 ;
        RECT 462.120000 515.540000 463.320000 516.020000 ;
        RECT 417.120000 515.540000 418.320000 516.020000 ;
        RECT 417.120000 493.780000 418.320000 494.260000 ;
        RECT 417.120000 488.340000 418.320000 488.820000 ;
        RECT 417.120000 482.900000 418.320000 483.380000 ;
        RECT 417.120000 499.220000 418.320000 499.700000 ;
        RECT 417.120000 504.660000 418.320000 505.140000 ;
        RECT 417.120000 510.100000 418.320000 510.580000 ;
        RECT 462.120000 493.780000 463.320000 494.260000 ;
        RECT 462.120000 488.340000 463.320000 488.820000 ;
        RECT 462.120000 482.900000 463.320000 483.380000 ;
        RECT 462.120000 504.660000 463.320000 505.140000 ;
        RECT 462.120000 499.220000 463.320000 499.700000 ;
        RECT 462.120000 510.100000 463.320000 510.580000 ;
        RECT 417.120000 520.980000 418.320000 521.460000 ;
        RECT 417.120000 526.420000 418.320000 526.900000 ;
        RECT 417.120000 531.860000 418.320000 532.340000 ;
        RECT 417.120000 537.300000 418.320000 537.780000 ;
        RECT 462.120000 520.980000 463.320000 521.460000 ;
        RECT 462.120000 526.420000 463.320000 526.900000 ;
        RECT 462.120000 531.860000 463.320000 532.340000 ;
        RECT 462.120000 537.300000 463.320000 537.780000 ;
        RECT 542.600000 515.540000 544.600000 516.020000 ;
        RECT 507.120000 515.540000 508.320000 516.020000 ;
        RECT 507.120000 488.340000 508.320000 488.820000 ;
        RECT 507.120000 482.900000 508.320000 483.380000 ;
        RECT 507.120000 493.780000 508.320000 494.260000 ;
        RECT 507.120000 499.220000 508.320000 499.700000 ;
        RECT 507.120000 504.660000 508.320000 505.140000 ;
        RECT 507.120000 510.100000 508.320000 510.580000 ;
        RECT 542.600000 493.780000 544.600000 494.260000 ;
        RECT 542.600000 488.340000 544.600000 488.820000 ;
        RECT 542.600000 482.900000 544.600000 483.380000 ;
        RECT 542.600000 510.100000 544.600000 510.580000 ;
        RECT 542.600000 504.660000 544.600000 505.140000 ;
        RECT 542.600000 499.220000 544.600000 499.700000 ;
        RECT 507.120000 526.420000 508.320000 526.900000 ;
        RECT 507.120000 520.980000 508.320000 521.460000 ;
        RECT 507.120000 531.860000 508.320000 532.340000 ;
        RECT 507.120000 537.300000 508.320000 537.780000 ;
        RECT 542.600000 531.860000 544.600000 532.340000 ;
        RECT 542.600000 526.420000 544.600000 526.900000 ;
        RECT 542.600000 520.980000 544.600000 521.460000 ;
        RECT 542.600000 537.300000 544.600000 537.780000 ;
      LAYER met4 ;
        RECT 507.120000 5.430000 508.320000 543.160000 ;
        RECT 462.120000 5.430000 463.320000 543.160000 ;
        RECT 417.120000 5.430000 418.320000 543.160000 ;
        RECT 372.120000 5.430000 373.320000 543.160000 ;
        RECT 327.120000 5.430000 328.320000 543.160000 ;
        RECT 282.120000 5.430000 283.320000 543.160000 ;
        RECT 237.120000 5.430000 238.320000 543.160000 ;
        RECT 192.120000 5.430000 193.320000 543.160000 ;
        RECT 147.120000 5.430000 148.320000 543.160000 ;
        RECT 102.120000 5.430000 103.320000 543.160000 ;
        RECT 57.120000 5.430000 58.320000 543.160000 ;
        RECT 12.120000 5.430000 13.320000 543.160000 ;
        RECT 542.600000 0.000000 544.600000 549.780000 ;
        RECT 5.560000 0.000000 7.560000 549.780000 ;
    END
# end of P/G power stripe data as pin

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 548.160000 544.160000 550.160000 546.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 544.160000 2.000000 546.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 548.160000 2.430000 550.160000 4.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 2.430000 2.000000 4.430000 ;
    END
    PORT
      LAYER met4 ;
        RECT 545.600000 547.780000 547.600000 549.780000 ;
    END
    PORT
      LAYER met4 ;
        RECT 545.600000 0.000000 547.600000 2.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.560000 547.780000 4.560000 549.780000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.560000 0.000000 4.560000 2.000000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 2.430000 550.160000 4.430000 ;
        RECT 0.000000 544.160000 550.160000 546.160000 ;
        RECT 2.560000 34.100000 4.560000 34.580000 ;
        RECT 9.955000 34.100000 11.320000 34.580000 ;
        RECT 55.120000 34.100000 56.320000 34.580000 ;
        RECT 2.560000 12.340000 4.560000 12.820000 ;
        RECT 9.955000 12.340000 11.320000 12.820000 ;
        RECT 2.560000 23.220000 4.560000 23.700000 ;
        RECT 9.955000 23.220000 11.320000 23.700000 ;
        RECT 2.560000 17.780000 4.560000 18.260000 ;
        RECT 9.955000 17.780000 11.320000 18.260000 ;
        RECT 2.560000 28.660000 4.560000 29.140000 ;
        RECT 9.955000 28.660000 11.320000 29.140000 ;
        RECT 55.120000 28.660000 56.320000 29.140000 ;
        RECT 55.120000 23.220000 56.320000 23.700000 ;
        RECT 55.120000 17.780000 56.320000 18.260000 ;
        RECT 55.120000 12.340000 56.320000 12.820000 ;
        RECT 2.560000 39.540000 4.560000 40.020000 ;
        RECT 9.955000 39.540000 11.320000 40.020000 ;
        RECT 2.560000 50.420000 4.560000 50.900000 ;
        RECT 9.955000 50.420000 11.320000 50.900000 ;
        RECT 2.560000 44.980000 4.560000 45.460000 ;
        RECT 9.955000 44.980000 11.320000 45.460000 ;
        RECT 2.560000 55.860000 4.560000 56.340000 ;
        RECT 9.955000 55.860000 11.320000 56.340000 ;
        RECT 2.560000 66.740000 4.560000 67.220000 ;
        RECT 9.955000 66.740000 11.320000 67.220000 ;
        RECT 2.560000 61.300000 4.560000 61.780000 ;
        RECT 9.955000 61.300000 11.320000 61.780000 ;
        RECT 55.120000 39.540000 56.320000 40.020000 ;
        RECT 55.120000 44.980000 56.320000 45.460000 ;
        RECT 55.120000 50.420000 56.320000 50.900000 ;
        RECT 55.120000 66.740000 56.320000 67.220000 ;
        RECT 55.120000 61.300000 56.320000 61.780000 ;
        RECT 55.120000 55.860000 56.320000 56.340000 ;
        RECT 100.120000 34.100000 101.320000 34.580000 ;
        RECT 100.120000 28.660000 101.320000 29.140000 ;
        RECT 100.120000 23.220000 101.320000 23.700000 ;
        RECT 100.120000 17.780000 101.320000 18.260000 ;
        RECT 100.120000 12.340000 101.320000 12.820000 ;
        RECT 100.120000 66.740000 101.320000 67.220000 ;
        RECT 100.120000 61.300000 101.320000 61.780000 ;
        RECT 100.120000 39.540000 101.320000 40.020000 ;
        RECT 100.120000 44.980000 101.320000 45.460000 ;
        RECT 100.120000 50.420000 101.320000 50.900000 ;
        RECT 100.120000 55.860000 101.320000 56.340000 ;
        RECT 2.560000 72.180000 4.560000 72.660000 ;
        RECT 9.955000 72.180000 11.320000 72.660000 ;
        RECT 2.560000 83.060000 4.560000 83.540000 ;
        RECT 9.955000 83.060000 11.320000 83.540000 ;
        RECT 2.560000 77.620000 4.560000 78.100000 ;
        RECT 9.955000 77.620000 11.320000 78.100000 ;
        RECT 2.560000 93.940000 4.560000 94.420000 ;
        RECT 9.955000 93.940000 11.320000 94.420000 ;
        RECT 2.560000 88.500000 4.560000 88.980000 ;
        RECT 9.955000 88.500000 11.320000 88.980000 ;
        RECT 2.560000 99.380000 4.560000 99.860000 ;
        RECT 9.955000 99.380000 11.320000 99.860000 ;
        RECT 55.120000 72.180000 56.320000 72.660000 ;
        RECT 55.120000 77.620000 56.320000 78.100000 ;
        RECT 55.120000 83.060000 56.320000 83.540000 ;
        RECT 55.120000 99.380000 56.320000 99.860000 ;
        RECT 55.120000 93.940000 56.320000 94.420000 ;
        RECT 55.120000 88.500000 56.320000 88.980000 ;
        RECT 2.560000 110.260000 4.560000 110.740000 ;
        RECT 9.955000 110.260000 11.320000 110.740000 ;
        RECT 2.560000 104.820000 4.560000 105.300000 ;
        RECT 9.955000 104.820000 11.320000 105.300000 ;
        RECT 2.560000 115.700000 4.560000 116.180000 ;
        RECT 9.955000 115.700000 11.320000 116.180000 ;
        RECT 2.560000 126.580000 4.560000 127.060000 ;
        RECT 9.955000 126.580000 11.320000 127.060000 ;
        RECT 2.560000 121.140000 4.560000 121.620000 ;
        RECT 9.955000 121.140000 11.320000 121.620000 ;
        RECT 2.560000 132.020000 4.560000 132.500000 ;
        RECT 9.955000 132.020000 11.320000 132.500000 ;
        RECT 55.120000 104.820000 56.320000 105.300000 ;
        RECT 55.120000 110.260000 56.320000 110.740000 ;
        RECT 55.120000 115.700000 56.320000 116.180000 ;
        RECT 55.120000 132.020000 56.320000 132.500000 ;
        RECT 55.120000 126.580000 56.320000 127.060000 ;
        RECT 55.120000 121.140000 56.320000 121.620000 ;
        RECT 100.120000 99.380000 101.320000 99.860000 ;
        RECT 100.120000 93.940000 101.320000 94.420000 ;
        RECT 100.120000 88.500000 101.320000 88.980000 ;
        RECT 100.120000 72.180000 101.320000 72.660000 ;
        RECT 100.120000 77.620000 101.320000 78.100000 ;
        RECT 100.120000 83.060000 101.320000 83.540000 ;
        RECT 100.120000 132.020000 101.320000 132.500000 ;
        RECT 100.120000 126.580000 101.320000 127.060000 ;
        RECT 100.120000 104.820000 101.320000 105.300000 ;
        RECT 100.120000 110.260000 101.320000 110.740000 ;
        RECT 100.120000 115.700000 101.320000 116.180000 ;
        RECT 100.120000 121.140000 101.320000 121.620000 ;
        RECT 190.120000 34.100000 191.320000 34.580000 ;
        RECT 145.120000 34.100000 146.320000 34.580000 ;
        RECT 145.120000 28.660000 146.320000 29.140000 ;
        RECT 145.120000 23.220000 146.320000 23.700000 ;
        RECT 145.120000 17.780000 146.320000 18.260000 ;
        RECT 145.120000 12.340000 146.320000 12.820000 ;
        RECT 190.120000 28.660000 191.320000 29.140000 ;
        RECT 190.120000 23.220000 191.320000 23.700000 ;
        RECT 190.120000 17.780000 191.320000 18.260000 ;
        RECT 190.120000 12.340000 191.320000 12.820000 ;
        RECT 145.120000 39.540000 146.320000 40.020000 ;
        RECT 145.120000 44.980000 146.320000 45.460000 ;
        RECT 145.120000 50.420000 146.320000 50.900000 ;
        RECT 145.120000 66.740000 146.320000 67.220000 ;
        RECT 145.120000 61.300000 146.320000 61.780000 ;
        RECT 145.120000 55.860000 146.320000 56.340000 ;
        RECT 190.120000 39.540000 191.320000 40.020000 ;
        RECT 190.120000 44.980000 191.320000 45.460000 ;
        RECT 190.120000 50.420000 191.320000 50.900000 ;
        RECT 190.120000 66.740000 191.320000 67.220000 ;
        RECT 190.120000 61.300000 191.320000 61.780000 ;
        RECT 190.120000 55.860000 191.320000 56.340000 ;
        RECT 235.120000 34.100000 236.320000 34.580000 ;
        RECT 235.120000 28.660000 236.320000 29.140000 ;
        RECT 235.120000 23.220000 236.320000 23.700000 ;
        RECT 235.120000 17.780000 236.320000 18.260000 ;
        RECT 235.120000 12.340000 236.320000 12.820000 ;
        RECT 235.120000 50.420000 236.320000 50.900000 ;
        RECT 235.120000 44.980000 236.320000 45.460000 ;
        RECT 235.120000 39.540000 236.320000 40.020000 ;
        RECT 235.120000 66.740000 236.320000 67.220000 ;
        RECT 235.120000 55.860000 236.320000 56.340000 ;
        RECT 235.120000 61.300000 236.320000 61.780000 ;
        RECT 145.120000 72.180000 146.320000 72.660000 ;
        RECT 145.120000 77.620000 146.320000 78.100000 ;
        RECT 145.120000 83.060000 146.320000 83.540000 ;
        RECT 145.120000 99.380000 146.320000 99.860000 ;
        RECT 145.120000 93.940000 146.320000 94.420000 ;
        RECT 145.120000 88.500000 146.320000 88.980000 ;
        RECT 190.120000 72.180000 191.320000 72.660000 ;
        RECT 190.120000 77.620000 191.320000 78.100000 ;
        RECT 190.120000 83.060000 191.320000 83.540000 ;
        RECT 190.120000 99.380000 191.320000 99.860000 ;
        RECT 190.120000 93.940000 191.320000 94.420000 ;
        RECT 190.120000 88.500000 191.320000 88.980000 ;
        RECT 145.120000 104.820000 146.320000 105.300000 ;
        RECT 145.120000 110.260000 146.320000 110.740000 ;
        RECT 145.120000 115.700000 146.320000 116.180000 ;
        RECT 145.120000 132.020000 146.320000 132.500000 ;
        RECT 145.120000 126.580000 146.320000 127.060000 ;
        RECT 145.120000 121.140000 146.320000 121.620000 ;
        RECT 190.120000 104.820000 191.320000 105.300000 ;
        RECT 190.120000 110.260000 191.320000 110.740000 ;
        RECT 190.120000 115.700000 191.320000 116.180000 ;
        RECT 190.120000 132.020000 191.320000 132.500000 ;
        RECT 190.120000 126.580000 191.320000 127.060000 ;
        RECT 190.120000 121.140000 191.320000 121.620000 ;
        RECT 235.120000 83.060000 236.320000 83.540000 ;
        RECT 235.120000 77.620000 236.320000 78.100000 ;
        RECT 235.120000 72.180000 236.320000 72.660000 ;
        RECT 235.120000 99.380000 236.320000 99.860000 ;
        RECT 235.120000 93.940000 236.320000 94.420000 ;
        RECT 235.120000 88.500000 236.320000 88.980000 ;
        RECT 235.120000 115.700000 236.320000 116.180000 ;
        RECT 235.120000 110.260000 236.320000 110.740000 ;
        RECT 235.120000 104.820000 236.320000 105.300000 ;
        RECT 235.120000 132.020000 236.320000 132.500000 ;
        RECT 235.120000 121.140000 236.320000 121.620000 ;
        RECT 235.120000 126.580000 236.320000 127.060000 ;
        RECT 2.560000 142.900000 4.560000 143.380000 ;
        RECT 9.955000 142.900000 11.320000 143.380000 ;
        RECT 2.560000 137.460000 4.560000 137.940000 ;
        RECT 9.955000 137.460000 11.320000 137.940000 ;
        RECT 2.560000 153.780000 4.560000 154.260000 ;
        RECT 9.955000 153.780000 11.320000 154.260000 ;
        RECT 2.560000 148.340000 4.560000 148.820000 ;
        RECT 9.955000 148.340000 11.320000 148.820000 ;
        RECT 2.560000 159.220000 4.560000 159.700000 ;
        RECT 9.955000 159.220000 11.320000 159.700000 ;
        RECT 2.560000 170.100000 4.560000 170.580000 ;
        RECT 9.955000 170.100000 11.320000 170.580000 ;
        RECT 2.560000 164.660000 4.560000 165.140000 ;
        RECT 9.955000 164.660000 11.320000 165.140000 ;
        RECT 55.120000 137.460000 56.320000 137.940000 ;
        RECT 55.120000 142.900000 56.320000 143.380000 ;
        RECT 55.120000 148.340000 56.320000 148.820000 ;
        RECT 55.120000 153.780000 56.320000 154.260000 ;
        RECT 55.120000 170.100000 56.320000 170.580000 ;
        RECT 55.120000 164.660000 56.320000 165.140000 ;
        RECT 55.120000 159.220000 56.320000 159.700000 ;
        RECT 2.560000 175.540000 4.560000 176.020000 ;
        RECT 9.955000 175.540000 11.320000 176.020000 ;
        RECT 2.560000 186.420000 4.560000 186.900000 ;
        RECT 9.955000 186.420000 11.320000 186.900000 ;
        RECT 2.560000 180.980000 4.560000 181.460000 ;
        RECT 9.955000 180.980000 11.320000 181.460000 ;
        RECT 2.560000 197.300000 4.560000 197.780000 ;
        RECT 9.955000 197.300000 11.320000 197.780000 ;
        RECT 2.560000 191.860000 4.560000 192.340000 ;
        RECT 9.955000 191.860000 11.320000 192.340000 ;
        RECT 2.560000 202.740000 4.560000 203.220000 ;
        RECT 9.955000 202.740000 11.320000 203.220000 ;
        RECT 55.120000 175.540000 56.320000 176.020000 ;
        RECT 55.120000 180.980000 56.320000 181.460000 ;
        RECT 55.120000 186.420000 56.320000 186.900000 ;
        RECT 55.120000 202.740000 56.320000 203.220000 ;
        RECT 55.120000 197.300000 56.320000 197.780000 ;
        RECT 55.120000 191.860000 56.320000 192.340000 ;
        RECT 100.120000 170.100000 101.320000 170.580000 ;
        RECT 100.120000 164.660000 101.320000 165.140000 ;
        RECT 100.120000 159.220000 101.320000 159.700000 ;
        RECT 100.120000 137.460000 101.320000 137.940000 ;
        RECT 100.120000 142.900000 101.320000 143.380000 ;
        RECT 100.120000 148.340000 101.320000 148.820000 ;
        RECT 100.120000 153.780000 101.320000 154.260000 ;
        RECT 100.120000 202.740000 101.320000 203.220000 ;
        RECT 100.120000 197.300000 101.320000 197.780000 ;
        RECT 100.120000 191.860000 101.320000 192.340000 ;
        RECT 100.120000 175.540000 101.320000 176.020000 ;
        RECT 100.120000 180.980000 101.320000 181.460000 ;
        RECT 100.120000 186.420000 101.320000 186.900000 ;
        RECT 2.560000 213.620000 4.560000 214.100000 ;
        RECT 9.955000 213.620000 11.320000 214.100000 ;
        RECT 2.560000 208.180000 4.560000 208.660000 ;
        RECT 9.955000 208.180000 11.320000 208.660000 ;
        RECT 2.560000 219.060000 4.560000 219.540000 ;
        RECT 9.955000 219.060000 11.320000 219.540000 ;
        RECT 2.560000 229.940000 4.560000 230.420000 ;
        RECT 9.955000 229.940000 11.320000 230.420000 ;
        RECT 2.560000 224.500000 4.560000 224.980000 ;
        RECT 9.955000 224.500000 11.320000 224.980000 ;
        RECT 2.560000 235.380000 4.560000 235.860000 ;
        RECT 9.955000 235.380000 11.320000 235.860000 ;
        RECT 55.120000 208.180000 56.320000 208.660000 ;
        RECT 55.120000 213.620000 56.320000 214.100000 ;
        RECT 55.120000 219.060000 56.320000 219.540000 ;
        RECT 55.120000 235.380000 56.320000 235.860000 ;
        RECT 55.120000 229.940000 56.320000 230.420000 ;
        RECT 55.120000 224.500000 56.320000 224.980000 ;
        RECT 2.560000 246.260000 4.560000 246.740000 ;
        RECT 9.955000 246.260000 11.320000 246.740000 ;
        RECT 2.560000 240.820000 4.560000 241.300000 ;
        RECT 9.955000 240.820000 11.320000 241.300000 ;
        RECT 2.560000 257.140000 4.560000 257.620000 ;
        RECT 9.955000 257.140000 11.320000 257.620000 ;
        RECT 2.560000 251.700000 4.560000 252.180000 ;
        RECT 9.955000 251.700000 11.320000 252.180000 ;
        RECT 2.560000 262.580000 4.560000 263.060000 ;
        RECT 9.955000 262.580000 11.320000 263.060000 ;
        RECT 2.560000 273.460000 4.560000 273.940000 ;
        RECT 9.955000 273.460000 11.320000 273.940000 ;
        RECT 2.560000 268.020000 4.560000 268.500000 ;
        RECT 9.955000 268.020000 11.320000 268.500000 ;
        RECT 55.120000 240.820000 56.320000 241.300000 ;
        RECT 55.120000 246.260000 56.320000 246.740000 ;
        RECT 55.120000 251.700000 56.320000 252.180000 ;
        RECT 55.120000 257.140000 56.320000 257.620000 ;
        RECT 55.120000 273.460000 56.320000 273.940000 ;
        RECT 55.120000 268.020000 56.320000 268.500000 ;
        RECT 55.120000 262.580000 56.320000 263.060000 ;
        RECT 100.120000 235.380000 101.320000 235.860000 ;
        RECT 100.120000 229.940000 101.320000 230.420000 ;
        RECT 100.120000 208.180000 101.320000 208.660000 ;
        RECT 100.120000 213.620000 101.320000 214.100000 ;
        RECT 100.120000 219.060000 101.320000 219.540000 ;
        RECT 100.120000 224.500000 101.320000 224.980000 ;
        RECT 100.120000 273.460000 101.320000 273.940000 ;
        RECT 100.120000 268.020000 101.320000 268.500000 ;
        RECT 100.120000 262.580000 101.320000 263.060000 ;
        RECT 100.120000 240.820000 101.320000 241.300000 ;
        RECT 100.120000 246.260000 101.320000 246.740000 ;
        RECT 100.120000 251.700000 101.320000 252.180000 ;
        RECT 100.120000 257.140000 101.320000 257.620000 ;
        RECT 145.120000 137.460000 146.320000 137.940000 ;
        RECT 145.120000 142.900000 146.320000 143.380000 ;
        RECT 145.120000 148.340000 146.320000 148.820000 ;
        RECT 145.120000 153.780000 146.320000 154.260000 ;
        RECT 145.120000 170.100000 146.320000 170.580000 ;
        RECT 145.120000 164.660000 146.320000 165.140000 ;
        RECT 145.120000 159.220000 146.320000 159.700000 ;
        RECT 190.120000 137.460000 191.320000 137.940000 ;
        RECT 190.120000 142.900000 191.320000 143.380000 ;
        RECT 190.120000 148.340000 191.320000 148.820000 ;
        RECT 190.120000 153.780000 191.320000 154.260000 ;
        RECT 190.120000 170.100000 191.320000 170.580000 ;
        RECT 190.120000 164.660000 191.320000 165.140000 ;
        RECT 190.120000 159.220000 191.320000 159.700000 ;
        RECT 145.120000 175.540000 146.320000 176.020000 ;
        RECT 145.120000 180.980000 146.320000 181.460000 ;
        RECT 145.120000 186.420000 146.320000 186.900000 ;
        RECT 145.120000 202.740000 146.320000 203.220000 ;
        RECT 145.120000 197.300000 146.320000 197.780000 ;
        RECT 145.120000 191.860000 146.320000 192.340000 ;
        RECT 190.120000 175.540000 191.320000 176.020000 ;
        RECT 190.120000 180.980000 191.320000 181.460000 ;
        RECT 190.120000 186.420000 191.320000 186.900000 ;
        RECT 190.120000 202.740000 191.320000 203.220000 ;
        RECT 190.120000 197.300000 191.320000 197.780000 ;
        RECT 190.120000 191.860000 191.320000 192.340000 ;
        RECT 235.120000 153.780000 236.320000 154.260000 ;
        RECT 235.120000 148.340000 236.320000 148.820000 ;
        RECT 235.120000 142.900000 236.320000 143.380000 ;
        RECT 235.120000 137.460000 236.320000 137.940000 ;
        RECT 235.120000 170.100000 236.320000 170.580000 ;
        RECT 235.120000 164.660000 236.320000 165.140000 ;
        RECT 235.120000 159.220000 236.320000 159.700000 ;
        RECT 235.120000 186.420000 236.320000 186.900000 ;
        RECT 235.120000 180.980000 236.320000 181.460000 ;
        RECT 235.120000 175.540000 236.320000 176.020000 ;
        RECT 235.120000 202.740000 236.320000 203.220000 ;
        RECT 235.120000 197.300000 236.320000 197.780000 ;
        RECT 235.120000 191.860000 236.320000 192.340000 ;
        RECT 145.120000 208.180000 146.320000 208.660000 ;
        RECT 145.120000 213.620000 146.320000 214.100000 ;
        RECT 145.120000 219.060000 146.320000 219.540000 ;
        RECT 145.120000 235.380000 146.320000 235.860000 ;
        RECT 145.120000 229.940000 146.320000 230.420000 ;
        RECT 145.120000 224.500000 146.320000 224.980000 ;
        RECT 190.120000 208.180000 191.320000 208.660000 ;
        RECT 190.120000 213.620000 191.320000 214.100000 ;
        RECT 190.120000 219.060000 191.320000 219.540000 ;
        RECT 190.120000 235.380000 191.320000 235.860000 ;
        RECT 190.120000 229.940000 191.320000 230.420000 ;
        RECT 190.120000 224.500000 191.320000 224.980000 ;
        RECT 145.120000 240.820000 146.320000 241.300000 ;
        RECT 145.120000 246.260000 146.320000 246.740000 ;
        RECT 145.120000 251.700000 146.320000 252.180000 ;
        RECT 145.120000 257.140000 146.320000 257.620000 ;
        RECT 145.120000 273.460000 146.320000 273.940000 ;
        RECT 145.120000 268.020000 146.320000 268.500000 ;
        RECT 145.120000 262.580000 146.320000 263.060000 ;
        RECT 190.120000 240.820000 191.320000 241.300000 ;
        RECT 190.120000 246.260000 191.320000 246.740000 ;
        RECT 190.120000 251.700000 191.320000 252.180000 ;
        RECT 190.120000 257.140000 191.320000 257.620000 ;
        RECT 190.120000 273.460000 191.320000 273.940000 ;
        RECT 190.120000 268.020000 191.320000 268.500000 ;
        RECT 190.120000 262.580000 191.320000 263.060000 ;
        RECT 235.120000 219.060000 236.320000 219.540000 ;
        RECT 235.120000 213.620000 236.320000 214.100000 ;
        RECT 235.120000 208.180000 236.320000 208.660000 ;
        RECT 235.120000 235.380000 236.320000 235.860000 ;
        RECT 235.120000 224.500000 236.320000 224.980000 ;
        RECT 235.120000 229.940000 236.320000 230.420000 ;
        RECT 235.120000 257.140000 236.320000 257.620000 ;
        RECT 235.120000 251.700000 236.320000 252.180000 ;
        RECT 235.120000 246.260000 236.320000 246.740000 ;
        RECT 235.120000 240.820000 236.320000 241.300000 ;
        RECT 235.120000 273.460000 236.320000 273.940000 ;
        RECT 235.120000 268.020000 236.320000 268.500000 ;
        RECT 235.120000 262.580000 236.320000 263.060000 ;
        RECT 325.120000 34.100000 326.320000 34.580000 ;
        RECT 280.120000 34.100000 281.320000 34.580000 ;
        RECT 280.120000 28.660000 281.320000 29.140000 ;
        RECT 280.120000 23.220000 281.320000 23.700000 ;
        RECT 280.120000 17.780000 281.320000 18.260000 ;
        RECT 280.120000 12.340000 281.320000 12.820000 ;
        RECT 325.120000 28.660000 326.320000 29.140000 ;
        RECT 325.120000 23.220000 326.320000 23.700000 ;
        RECT 325.120000 17.780000 326.320000 18.260000 ;
        RECT 325.120000 12.340000 326.320000 12.820000 ;
        RECT 280.120000 39.540000 281.320000 40.020000 ;
        RECT 280.120000 44.980000 281.320000 45.460000 ;
        RECT 280.120000 50.420000 281.320000 50.900000 ;
        RECT 280.120000 66.740000 281.320000 67.220000 ;
        RECT 280.120000 61.300000 281.320000 61.780000 ;
        RECT 280.120000 55.860000 281.320000 56.340000 ;
        RECT 325.120000 39.540000 326.320000 40.020000 ;
        RECT 325.120000 44.980000 326.320000 45.460000 ;
        RECT 325.120000 50.420000 326.320000 50.900000 ;
        RECT 325.120000 66.740000 326.320000 67.220000 ;
        RECT 325.120000 61.300000 326.320000 61.780000 ;
        RECT 325.120000 55.860000 326.320000 56.340000 ;
        RECT 370.120000 34.100000 371.320000 34.580000 ;
        RECT 370.120000 28.660000 371.320000 29.140000 ;
        RECT 370.120000 23.220000 371.320000 23.700000 ;
        RECT 370.120000 17.780000 371.320000 18.260000 ;
        RECT 370.120000 12.340000 371.320000 12.820000 ;
        RECT 370.120000 50.420000 371.320000 50.900000 ;
        RECT 370.120000 44.980000 371.320000 45.460000 ;
        RECT 370.120000 39.540000 371.320000 40.020000 ;
        RECT 370.120000 66.740000 371.320000 67.220000 ;
        RECT 370.120000 55.860000 371.320000 56.340000 ;
        RECT 370.120000 61.300000 371.320000 61.780000 ;
        RECT 280.120000 72.180000 281.320000 72.660000 ;
        RECT 280.120000 77.620000 281.320000 78.100000 ;
        RECT 280.120000 83.060000 281.320000 83.540000 ;
        RECT 280.120000 99.380000 281.320000 99.860000 ;
        RECT 280.120000 93.940000 281.320000 94.420000 ;
        RECT 280.120000 88.500000 281.320000 88.980000 ;
        RECT 325.120000 72.180000 326.320000 72.660000 ;
        RECT 325.120000 77.620000 326.320000 78.100000 ;
        RECT 325.120000 83.060000 326.320000 83.540000 ;
        RECT 325.120000 99.380000 326.320000 99.860000 ;
        RECT 325.120000 93.940000 326.320000 94.420000 ;
        RECT 325.120000 88.500000 326.320000 88.980000 ;
        RECT 280.120000 104.820000 281.320000 105.300000 ;
        RECT 280.120000 110.260000 281.320000 110.740000 ;
        RECT 280.120000 115.700000 281.320000 116.180000 ;
        RECT 280.120000 132.020000 281.320000 132.500000 ;
        RECT 280.120000 126.580000 281.320000 127.060000 ;
        RECT 280.120000 121.140000 281.320000 121.620000 ;
        RECT 325.120000 104.820000 326.320000 105.300000 ;
        RECT 325.120000 110.260000 326.320000 110.740000 ;
        RECT 325.120000 115.700000 326.320000 116.180000 ;
        RECT 325.120000 132.020000 326.320000 132.500000 ;
        RECT 325.120000 126.580000 326.320000 127.060000 ;
        RECT 325.120000 121.140000 326.320000 121.620000 ;
        RECT 370.120000 83.060000 371.320000 83.540000 ;
        RECT 370.120000 77.620000 371.320000 78.100000 ;
        RECT 370.120000 72.180000 371.320000 72.660000 ;
        RECT 370.120000 99.380000 371.320000 99.860000 ;
        RECT 370.120000 93.940000 371.320000 94.420000 ;
        RECT 370.120000 88.500000 371.320000 88.980000 ;
        RECT 370.120000 115.700000 371.320000 116.180000 ;
        RECT 370.120000 110.260000 371.320000 110.740000 ;
        RECT 370.120000 104.820000 371.320000 105.300000 ;
        RECT 370.120000 132.020000 371.320000 132.500000 ;
        RECT 370.120000 121.140000 371.320000 121.620000 ;
        RECT 370.120000 126.580000 371.320000 127.060000 ;
        RECT 460.120000 34.100000 461.320000 34.580000 ;
        RECT 415.120000 34.100000 416.320000 34.580000 ;
        RECT 415.120000 28.660000 416.320000 29.140000 ;
        RECT 415.120000 23.220000 416.320000 23.700000 ;
        RECT 415.120000 17.780000 416.320000 18.260000 ;
        RECT 415.120000 12.340000 416.320000 12.820000 ;
        RECT 460.120000 28.660000 461.320000 29.140000 ;
        RECT 460.120000 23.220000 461.320000 23.700000 ;
        RECT 460.120000 17.780000 461.320000 18.260000 ;
        RECT 460.120000 12.340000 461.320000 12.820000 ;
        RECT 415.120000 39.540000 416.320000 40.020000 ;
        RECT 415.120000 44.980000 416.320000 45.460000 ;
        RECT 415.120000 50.420000 416.320000 50.900000 ;
        RECT 415.120000 66.740000 416.320000 67.220000 ;
        RECT 415.120000 61.300000 416.320000 61.780000 ;
        RECT 415.120000 55.860000 416.320000 56.340000 ;
        RECT 460.120000 39.540000 461.320000 40.020000 ;
        RECT 460.120000 44.980000 461.320000 45.460000 ;
        RECT 460.120000 50.420000 461.320000 50.900000 ;
        RECT 460.120000 66.740000 461.320000 67.220000 ;
        RECT 460.120000 61.300000 461.320000 61.780000 ;
        RECT 460.120000 55.860000 461.320000 56.340000 ;
        RECT 545.600000 34.100000 547.600000 34.580000 ;
        RECT 505.120000 34.100000 506.320000 34.580000 ;
        RECT 505.120000 12.340000 506.320000 12.820000 ;
        RECT 505.120000 17.780000 506.320000 18.260000 ;
        RECT 505.120000 23.220000 506.320000 23.700000 ;
        RECT 505.120000 28.660000 506.320000 29.140000 ;
        RECT 545.600000 12.340000 547.600000 12.820000 ;
        RECT 545.600000 28.660000 547.600000 29.140000 ;
        RECT 545.600000 23.220000 547.600000 23.700000 ;
        RECT 545.600000 17.780000 547.600000 18.260000 ;
        RECT 505.120000 50.420000 506.320000 50.900000 ;
        RECT 505.120000 44.980000 506.320000 45.460000 ;
        RECT 505.120000 39.540000 506.320000 40.020000 ;
        RECT 505.120000 66.740000 506.320000 67.220000 ;
        RECT 505.120000 55.860000 506.320000 56.340000 ;
        RECT 505.120000 61.300000 506.320000 61.780000 ;
        RECT 545.600000 50.420000 547.600000 50.900000 ;
        RECT 545.600000 39.540000 547.600000 40.020000 ;
        RECT 545.600000 44.980000 547.600000 45.460000 ;
        RECT 545.600000 66.740000 547.600000 67.220000 ;
        RECT 545.600000 61.300000 547.600000 61.780000 ;
        RECT 545.600000 55.860000 547.600000 56.340000 ;
        RECT 415.120000 72.180000 416.320000 72.660000 ;
        RECT 415.120000 77.620000 416.320000 78.100000 ;
        RECT 415.120000 83.060000 416.320000 83.540000 ;
        RECT 415.120000 99.380000 416.320000 99.860000 ;
        RECT 415.120000 93.940000 416.320000 94.420000 ;
        RECT 415.120000 88.500000 416.320000 88.980000 ;
        RECT 460.120000 72.180000 461.320000 72.660000 ;
        RECT 460.120000 77.620000 461.320000 78.100000 ;
        RECT 460.120000 83.060000 461.320000 83.540000 ;
        RECT 460.120000 99.380000 461.320000 99.860000 ;
        RECT 460.120000 93.940000 461.320000 94.420000 ;
        RECT 460.120000 88.500000 461.320000 88.980000 ;
        RECT 415.120000 104.820000 416.320000 105.300000 ;
        RECT 415.120000 110.260000 416.320000 110.740000 ;
        RECT 415.120000 115.700000 416.320000 116.180000 ;
        RECT 415.120000 132.020000 416.320000 132.500000 ;
        RECT 415.120000 126.580000 416.320000 127.060000 ;
        RECT 415.120000 121.140000 416.320000 121.620000 ;
        RECT 460.120000 104.820000 461.320000 105.300000 ;
        RECT 460.120000 110.260000 461.320000 110.740000 ;
        RECT 460.120000 115.700000 461.320000 116.180000 ;
        RECT 460.120000 132.020000 461.320000 132.500000 ;
        RECT 460.120000 126.580000 461.320000 127.060000 ;
        RECT 460.120000 121.140000 461.320000 121.620000 ;
        RECT 505.120000 83.060000 506.320000 83.540000 ;
        RECT 505.120000 77.620000 506.320000 78.100000 ;
        RECT 505.120000 72.180000 506.320000 72.660000 ;
        RECT 505.120000 99.380000 506.320000 99.860000 ;
        RECT 505.120000 93.940000 506.320000 94.420000 ;
        RECT 505.120000 88.500000 506.320000 88.980000 ;
        RECT 545.600000 83.060000 547.600000 83.540000 ;
        RECT 545.600000 77.620000 547.600000 78.100000 ;
        RECT 545.600000 72.180000 547.600000 72.660000 ;
        RECT 545.600000 99.380000 547.600000 99.860000 ;
        RECT 545.600000 93.940000 547.600000 94.420000 ;
        RECT 545.600000 88.500000 547.600000 88.980000 ;
        RECT 505.120000 115.700000 506.320000 116.180000 ;
        RECT 505.120000 110.260000 506.320000 110.740000 ;
        RECT 505.120000 104.820000 506.320000 105.300000 ;
        RECT 505.120000 132.020000 506.320000 132.500000 ;
        RECT 505.120000 121.140000 506.320000 121.620000 ;
        RECT 505.120000 126.580000 506.320000 127.060000 ;
        RECT 545.600000 115.700000 547.600000 116.180000 ;
        RECT 545.600000 104.820000 547.600000 105.300000 ;
        RECT 545.600000 110.260000 547.600000 110.740000 ;
        RECT 545.600000 132.020000 547.600000 132.500000 ;
        RECT 545.600000 126.580000 547.600000 127.060000 ;
        RECT 545.600000 121.140000 547.600000 121.620000 ;
        RECT 280.120000 137.460000 281.320000 137.940000 ;
        RECT 280.120000 142.900000 281.320000 143.380000 ;
        RECT 280.120000 148.340000 281.320000 148.820000 ;
        RECT 280.120000 153.780000 281.320000 154.260000 ;
        RECT 280.120000 170.100000 281.320000 170.580000 ;
        RECT 280.120000 164.660000 281.320000 165.140000 ;
        RECT 280.120000 159.220000 281.320000 159.700000 ;
        RECT 325.120000 137.460000 326.320000 137.940000 ;
        RECT 325.120000 142.900000 326.320000 143.380000 ;
        RECT 325.120000 148.340000 326.320000 148.820000 ;
        RECT 325.120000 153.780000 326.320000 154.260000 ;
        RECT 325.120000 170.100000 326.320000 170.580000 ;
        RECT 325.120000 164.660000 326.320000 165.140000 ;
        RECT 325.120000 159.220000 326.320000 159.700000 ;
        RECT 280.120000 175.540000 281.320000 176.020000 ;
        RECT 280.120000 180.980000 281.320000 181.460000 ;
        RECT 280.120000 186.420000 281.320000 186.900000 ;
        RECT 280.120000 202.740000 281.320000 203.220000 ;
        RECT 280.120000 197.300000 281.320000 197.780000 ;
        RECT 280.120000 191.860000 281.320000 192.340000 ;
        RECT 325.120000 175.540000 326.320000 176.020000 ;
        RECT 325.120000 180.980000 326.320000 181.460000 ;
        RECT 325.120000 186.420000 326.320000 186.900000 ;
        RECT 325.120000 202.740000 326.320000 203.220000 ;
        RECT 325.120000 197.300000 326.320000 197.780000 ;
        RECT 325.120000 191.860000 326.320000 192.340000 ;
        RECT 370.120000 153.780000 371.320000 154.260000 ;
        RECT 370.120000 148.340000 371.320000 148.820000 ;
        RECT 370.120000 142.900000 371.320000 143.380000 ;
        RECT 370.120000 137.460000 371.320000 137.940000 ;
        RECT 370.120000 170.100000 371.320000 170.580000 ;
        RECT 370.120000 164.660000 371.320000 165.140000 ;
        RECT 370.120000 159.220000 371.320000 159.700000 ;
        RECT 370.120000 186.420000 371.320000 186.900000 ;
        RECT 370.120000 180.980000 371.320000 181.460000 ;
        RECT 370.120000 175.540000 371.320000 176.020000 ;
        RECT 370.120000 202.740000 371.320000 203.220000 ;
        RECT 370.120000 197.300000 371.320000 197.780000 ;
        RECT 370.120000 191.860000 371.320000 192.340000 ;
        RECT 280.120000 208.180000 281.320000 208.660000 ;
        RECT 280.120000 213.620000 281.320000 214.100000 ;
        RECT 280.120000 219.060000 281.320000 219.540000 ;
        RECT 280.120000 235.380000 281.320000 235.860000 ;
        RECT 280.120000 229.940000 281.320000 230.420000 ;
        RECT 280.120000 224.500000 281.320000 224.980000 ;
        RECT 325.120000 208.180000 326.320000 208.660000 ;
        RECT 325.120000 213.620000 326.320000 214.100000 ;
        RECT 325.120000 219.060000 326.320000 219.540000 ;
        RECT 325.120000 235.380000 326.320000 235.860000 ;
        RECT 325.120000 229.940000 326.320000 230.420000 ;
        RECT 325.120000 224.500000 326.320000 224.980000 ;
        RECT 280.120000 240.820000 281.320000 241.300000 ;
        RECT 280.120000 246.260000 281.320000 246.740000 ;
        RECT 280.120000 251.700000 281.320000 252.180000 ;
        RECT 280.120000 257.140000 281.320000 257.620000 ;
        RECT 280.120000 273.460000 281.320000 273.940000 ;
        RECT 280.120000 268.020000 281.320000 268.500000 ;
        RECT 280.120000 262.580000 281.320000 263.060000 ;
        RECT 325.120000 240.820000 326.320000 241.300000 ;
        RECT 325.120000 246.260000 326.320000 246.740000 ;
        RECT 325.120000 251.700000 326.320000 252.180000 ;
        RECT 325.120000 257.140000 326.320000 257.620000 ;
        RECT 325.120000 273.460000 326.320000 273.940000 ;
        RECT 325.120000 268.020000 326.320000 268.500000 ;
        RECT 325.120000 262.580000 326.320000 263.060000 ;
        RECT 370.120000 219.060000 371.320000 219.540000 ;
        RECT 370.120000 213.620000 371.320000 214.100000 ;
        RECT 370.120000 208.180000 371.320000 208.660000 ;
        RECT 370.120000 235.380000 371.320000 235.860000 ;
        RECT 370.120000 224.500000 371.320000 224.980000 ;
        RECT 370.120000 229.940000 371.320000 230.420000 ;
        RECT 370.120000 257.140000 371.320000 257.620000 ;
        RECT 370.120000 251.700000 371.320000 252.180000 ;
        RECT 370.120000 246.260000 371.320000 246.740000 ;
        RECT 370.120000 240.820000 371.320000 241.300000 ;
        RECT 370.120000 273.460000 371.320000 273.940000 ;
        RECT 370.120000 268.020000 371.320000 268.500000 ;
        RECT 370.120000 262.580000 371.320000 263.060000 ;
        RECT 415.120000 137.460000 416.320000 137.940000 ;
        RECT 415.120000 142.900000 416.320000 143.380000 ;
        RECT 415.120000 148.340000 416.320000 148.820000 ;
        RECT 415.120000 153.780000 416.320000 154.260000 ;
        RECT 415.120000 170.100000 416.320000 170.580000 ;
        RECT 415.120000 164.660000 416.320000 165.140000 ;
        RECT 415.120000 159.220000 416.320000 159.700000 ;
        RECT 460.120000 137.460000 461.320000 137.940000 ;
        RECT 460.120000 142.900000 461.320000 143.380000 ;
        RECT 460.120000 148.340000 461.320000 148.820000 ;
        RECT 460.120000 153.780000 461.320000 154.260000 ;
        RECT 460.120000 170.100000 461.320000 170.580000 ;
        RECT 460.120000 164.660000 461.320000 165.140000 ;
        RECT 460.120000 159.220000 461.320000 159.700000 ;
        RECT 415.120000 175.540000 416.320000 176.020000 ;
        RECT 415.120000 180.980000 416.320000 181.460000 ;
        RECT 415.120000 186.420000 416.320000 186.900000 ;
        RECT 415.120000 202.740000 416.320000 203.220000 ;
        RECT 415.120000 197.300000 416.320000 197.780000 ;
        RECT 415.120000 191.860000 416.320000 192.340000 ;
        RECT 460.120000 175.540000 461.320000 176.020000 ;
        RECT 460.120000 180.980000 461.320000 181.460000 ;
        RECT 460.120000 186.420000 461.320000 186.900000 ;
        RECT 460.120000 202.740000 461.320000 203.220000 ;
        RECT 460.120000 197.300000 461.320000 197.780000 ;
        RECT 460.120000 191.860000 461.320000 192.340000 ;
        RECT 505.120000 153.780000 506.320000 154.260000 ;
        RECT 505.120000 148.340000 506.320000 148.820000 ;
        RECT 505.120000 142.900000 506.320000 143.380000 ;
        RECT 505.120000 137.460000 506.320000 137.940000 ;
        RECT 505.120000 170.100000 506.320000 170.580000 ;
        RECT 505.120000 164.660000 506.320000 165.140000 ;
        RECT 505.120000 159.220000 506.320000 159.700000 ;
        RECT 545.600000 153.780000 547.600000 154.260000 ;
        RECT 545.600000 148.340000 547.600000 148.820000 ;
        RECT 545.600000 137.460000 547.600000 137.940000 ;
        RECT 545.600000 142.900000 547.600000 143.380000 ;
        RECT 545.600000 170.100000 547.600000 170.580000 ;
        RECT 545.600000 164.660000 547.600000 165.140000 ;
        RECT 545.600000 159.220000 547.600000 159.700000 ;
        RECT 505.120000 186.420000 506.320000 186.900000 ;
        RECT 505.120000 180.980000 506.320000 181.460000 ;
        RECT 505.120000 175.540000 506.320000 176.020000 ;
        RECT 505.120000 202.740000 506.320000 203.220000 ;
        RECT 505.120000 197.300000 506.320000 197.780000 ;
        RECT 505.120000 191.860000 506.320000 192.340000 ;
        RECT 545.600000 186.420000 547.600000 186.900000 ;
        RECT 545.600000 180.980000 547.600000 181.460000 ;
        RECT 545.600000 175.540000 547.600000 176.020000 ;
        RECT 545.600000 202.740000 547.600000 203.220000 ;
        RECT 545.600000 197.300000 547.600000 197.780000 ;
        RECT 545.600000 191.860000 547.600000 192.340000 ;
        RECT 415.120000 208.180000 416.320000 208.660000 ;
        RECT 415.120000 213.620000 416.320000 214.100000 ;
        RECT 415.120000 219.060000 416.320000 219.540000 ;
        RECT 415.120000 235.380000 416.320000 235.860000 ;
        RECT 415.120000 229.940000 416.320000 230.420000 ;
        RECT 415.120000 224.500000 416.320000 224.980000 ;
        RECT 460.120000 208.180000 461.320000 208.660000 ;
        RECT 460.120000 213.620000 461.320000 214.100000 ;
        RECT 460.120000 219.060000 461.320000 219.540000 ;
        RECT 460.120000 235.380000 461.320000 235.860000 ;
        RECT 460.120000 229.940000 461.320000 230.420000 ;
        RECT 460.120000 224.500000 461.320000 224.980000 ;
        RECT 415.120000 240.820000 416.320000 241.300000 ;
        RECT 415.120000 246.260000 416.320000 246.740000 ;
        RECT 415.120000 251.700000 416.320000 252.180000 ;
        RECT 415.120000 257.140000 416.320000 257.620000 ;
        RECT 415.120000 273.460000 416.320000 273.940000 ;
        RECT 415.120000 268.020000 416.320000 268.500000 ;
        RECT 415.120000 262.580000 416.320000 263.060000 ;
        RECT 460.120000 240.820000 461.320000 241.300000 ;
        RECT 460.120000 246.260000 461.320000 246.740000 ;
        RECT 460.120000 251.700000 461.320000 252.180000 ;
        RECT 460.120000 257.140000 461.320000 257.620000 ;
        RECT 460.120000 273.460000 461.320000 273.940000 ;
        RECT 460.120000 268.020000 461.320000 268.500000 ;
        RECT 460.120000 262.580000 461.320000 263.060000 ;
        RECT 505.120000 219.060000 506.320000 219.540000 ;
        RECT 505.120000 213.620000 506.320000 214.100000 ;
        RECT 505.120000 208.180000 506.320000 208.660000 ;
        RECT 505.120000 235.380000 506.320000 235.860000 ;
        RECT 505.120000 224.500000 506.320000 224.980000 ;
        RECT 505.120000 229.940000 506.320000 230.420000 ;
        RECT 545.600000 219.060000 547.600000 219.540000 ;
        RECT 545.600000 208.180000 547.600000 208.660000 ;
        RECT 545.600000 213.620000 547.600000 214.100000 ;
        RECT 545.600000 235.380000 547.600000 235.860000 ;
        RECT 545.600000 229.940000 547.600000 230.420000 ;
        RECT 545.600000 224.500000 547.600000 224.980000 ;
        RECT 505.120000 257.140000 506.320000 257.620000 ;
        RECT 505.120000 251.700000 506.320000 252.180000 ;
        RECT 505.120000 246.260000 506.320000 246.740000 ;
        RECT 505.120000 240.820000 506.320000 241.300000 ;
        RECT 505.120000 273.460000 506.320000 273.940000 ;
        RECT 505.120000 268.020000 506.320000 268.500000 ;
        RECT 505.120000 262.580000 506.320000 263.060000 ;
        RECT 545.600000 257.140000 547.600000 257.620000 ;
        RECT 545.600000 251.700000 547.600000 252.180000 ;
        RECT 545.600000 240.820000 547.600000 241.300000 ;
        RECT 545.600000 246.260000 547.600000 246.740000 ;
        RECT 545.600000 273.460000 547.600000 273.940000 ;
        RECT 545.600000 268.020000 547.600000 268.500000 ;
        RECT 545.600000 262.580000 547.600000 263.060000 ;
        RECT 2.560000 278.900000 4.560000 279.380000 ;
        RECT 9.955000 278.900000 11.320000 279.380000 ;
        RECT 2.560000 289.780000 4.560000 290.260000 ;
        RECT 9.955000 289.780000 11.320000 290.260000 ;
        RECT 2.560000 284.340000 4.560000 284.820000 ;
        RECT 9.955000 284.340000 11.320000 284.820000 ;
        RECT 2.560000 300.660000 4.560000 301.140000 ;
        RECT 9.955000 300.660000 11.320000 301.140000 ;
        RECT 2.560000 295.220000 4.560000 295.700000 ;
        RECT 9.955000 295.220000 11.320000 295.700000 ;
        RECT 2.560000 306.100000 4.560000 306.580000 ;
        RECT 9.955000 306.100000 11.320000 306.580000 ;
        RECT 55.120000 278.900000 56.320000 279.380000 ;
        RECT 55.120000 284.340000 56.320000 284.820000 ;
        RECT 55.120000 289.780000 56.320000 290.260000 ;
        RECT 55.120000 306.100000 56.320000 306.580000 ;
        RECT 55.120000 300.660000 56.320000 301.140000 ;
        RECT 55.120000 295.220000 56.320000 295.700000 ;
        RECT 2.560000 316.980000 4.560000 317.460000 ;
        RECT 9.955000 316.980000 11.320000 317.460000 ;
        RECT 2.560000 311.540000 4.560000 312.020000 ;
        RECT 9.955000 311.540000 11.320000 312.020000 ;
        RECT 2.560000 322.420000 4.560000 322.900000 ;
        RECT 9.955000 322.420000 11.320000 322.900000 ;
        RECT 2.560000 333.300000 4.560000 333.780000 ;
        RECT 9.955000 333.300000 11.320000 333.780000 ;
        RECT 2.560000 327.860000 4.560000 328.340000 ;
        RECT 9.955000 327.860000 11.320000 328.340000 ;
        RECT 2.560000 338.740000 4.560000 339.220000 ;
        RECT 9.955000 338.740000 11.320000 339.220000 ;
        RECT 55.120000 311.540000 56.320000 312.020000 ;
        RECT 55.120000 316.980000 56.320000 317.460000 ;
        RECT 55.120000 322.420000 56.320000 322.900000 ;
        RECT 55.120000 338.740000 56.320000 339.220000 ;
        RECT 55.120000 333.300000 56.320000 333.780000 ;
        RECT 55.120000 327.860000 56.320000 328.340000 ;
        RECT 100.120000 306.100000 101.320000 306.580000 ;
        RECT 100.120000 300.660000 101.320000 301.140000 ;
        RECT 100.120000 278.900000 101.320000 279.380000 ;
        RECT 100.120000 284.340000 101.320000 284.820000 ;
        RECT 100.120000 289.780000 101.320000 290.260000 ;
        RECT 100.120000 295.220000 101.320000 295.700000 ;
        RECT 100.120000 338.740000 101.320000 339.220000 ;
        RECT 100.120000 333.300000 101.320000 333.780000 ;
        RECT 100.120000 311.540000 101.320000 312.020000 ;
        RECT 100.120000 316.980000 101.320000 317.460000 ;
        RECT 100.120000 322.420000 101.320000 322.900000 ;
        RECT 100.120000 327.860000 101.320000 328.340000 ;
        RECT 2.560000 360.500000 4.560000 360.980000 ;
        RECT 9.955000 360.500000 11.320000 360.980000 ;
        RECT 2.560000 349.620000 4.560000 350.100000 ;
        RECT 9.955000 349.620000 11.320000 350.100000 ;
        RECT 2.560000 344.180000 4.560000 344.660000 ;
        RECT 9.955000 344.180000 11.320000 344.660000 ;
        RECT 2.560000 355.060000 4.560000 355.540000 ;
        RECT 9.955000 355.060000 11.320000 355.540000 ;
        RECT 2.560000 365.940000 4.560000 366.420000 ;
        RECT 9.955000 365.940000 11.320000 366.420000 ;
        RECT 2.560000 376.820000 4.560000 377.300000 ;
        RECT 9.955000 376.820000 11.320000 377.300000 ;
        RECT 2.560000 371.380000 4.560000 371.860000 ;
        RECT 9.955000 371.380000 11.320000 371.860000 ;
        RECT 55.120000 360.500000 56.320000 360.980000 ;
        RECT 55.120000 344.180000 56.320000 344.660000 ;
        RECT 55.120000 349.620000 56.320000 350.100000 ;
        RECT 55.120000 355.060000 56.320000 355.540000 ;
        RECT 55.120000 376.820000 56.320000 377.300000 ;
        RECT 55.120000 371.380000 56.320000 371.860000 ;
        RECT 55.120000 365.940000 56.320000 366.420000 ;
        RECT 2.560000 382.260000 4.560000 382.740000 ;
        RECT 9.955000 382.260000 11.320000 382.740000 ;
        RECT 2.560000 393.140000 4.560000 393.620000 ;
        RECT 9.955000 393.140000 11.320000 393.620000 ;
        RECT 2.560000 387.700000 4.560000 388.180000 ;
        RECT 9.955000 387.700000 11.320000 388.180000 ;
        RECT 2.560000 398.580000 4.560000 399.060000 ;
        RECT 9.955000 398.580000 11.320000 399.060000 ;
        RECT 2.560000 409.460000 4.560000 409.940000 ;
        RECT 9.955000 409.460000 11.320000 409.940000 ;
        RECT 2.560000 404.020000 4.560000 404.500000 ;
        RECT 9.955000 404.020000 11.320000 404.500000 ;
        RECT 55.120000 382.260000 56.320000 382.740000 ;
        RECT 55.120000 387.700000 56.320000 388.180000 ;
        RECT 55.120000 393.140000 56.320000 393.620000 ;
        RECT 55.120000 409.460000 56.320000 409.940000 ;
        RECT 55.120000 404.020000 56.320000 404.500000 ;
        RECT 55.120000 398.580000 56.320000 399.060000 ;
        RECT 100.120000 376.820000 101.320000 377.300000 ;
        RECT 100.120000 371.380000 101.320000 371.860000 ;
        RECT 100.120000 365.940000 101.320000 366.420000 ;
        RECT 100.120000 344.180000 101.320000 344.660000 ;
        RECT 100.120000 349.620000 101.320000 350.100000 ;
        RECT 100.120000 355.060000 101.320000 355.540000 ;
        RECT 100.120000 360.500000 101.320000 360.980000 ;
        RECT 100.120000 409.460000 101.320000 409.940000 ;
        RECT 100.120000 404.020000 101.320000 404.500000 ;
        RECT 100.120000 382.260000 101.320000 382.740000 ;
        RECT 100.120000 387.700000 101.320000 388.180000 ;
        RECT 100.120000 393.140000 101.320000 393.620000 ;
        RECT 100.120000 398.580000 101.320000 399.060000 ;
        RECT 145.120000 278.900000 146.320000 279.380000 ;
        RECT 145.120000 284.340000 146.320000 284.820000 ;
        RECT 145.120000 289.780000 146.320000 290.260000 ;
        RECT 145.120000 306.100000 146.320000 306.580000 ;
        RECT 145.120000 300.660000 146.320000 301.140000 ;
        RECT 145.120000 295.220000 146.320000 295.700000 ;
        RECT 190.120000 278.900000 191.320000 279.380000 ;
        RECT 190.120000 284.340000 191.320000 284.820000 ;
        RECT 190.120000 289.780000 191.320000 290.260000 ;
        RECT 190.120000 306.100000 191.320000 306.580000 ;
        RECT 190.120000 300.660000 191.320000 301.140000 ;
        RECT 190.120000 295.220000 191.320000 295.700000 ;
        RECT 145.120000 311.540000 146.320000 312.020000 ;
        RECT 145.120000 316.980000 146.320000 317.460000 ;
        RECT 145.120000 322.420000 146.320000 322.900000 ;
        RECT 145.120000 338.740000 146.320000 339.220000 ;
        RECT 145.120000 333.300000 146.320000 333.780000 ;
        RECT 145.120000 327.860000 146.320000 328.340000 ;
        RECT 190.120000 311.540000 191.320000 312.020000 ;
        RECT 190.120000 316.980000 191.320000 317.460000 ;
        RECT 190.120000 322.420000 191.320000 322.900000 ;
        RECT 190.120000 338.740000 191.320000 339.220000 ;
        RECT 190.120000 333.300000 191.320000 333.780000 ;
        RECT 190.120000 327.860000 191.320000 328.340000 ;
        RECT 235.120000 289.780000 236.320000 290.260000 ;
        RECT 235.120000 284.340000 236.320000 284.820000 ;
        RECT 235.120000 278.900000 236.320000 279.380000 ;
        RECT 235.120000 306.100000 236.320000 306.580000 ;
        RECT 235.120000 295.220000 236.320000 295.700000 ;
        RECT 235.120000 300.660000 236.320000 301.140000 ;
        RECT 235.120000 322.420000 236.320000 322.900000 ;
        RECT 235.120000 316.980000 236.320000 317.460000 ;
        RECT 235.120000 311.540000 236.320000 312.020000 ;
        RECT 235.120000 338.740000 236.320000 339.220000 ;
        RECT 235.120000 327.860000 236.320000 328.340000 ;
        RECT 235.120000 333.300000 236.320000 333.780000 ;
        RECT 145.120000 360.500000 146.320000 360.980000 ;
        RECT 145.120000 344.180000 146.320000 344.660000 ;
        RECT 145.120000 349.620000 146.320000 350.100000 ;
        RECT 145.120000 355.060000 146.320000 355.540000 ;
        RECT 145.120000 376.820000 146.320000 377.300000 ;
        RECT 145.120000 371.380000 146.320000 371.860000 ;
        RECT 145.120000 365.940000 146.320000 366.420000 ;
        RECT 190.120000 360.500000 191.320000 360.980000 ;
        RECT 190.120000 344.180000 191.320000 344.660000 ;
        RECT 190.120000 349.620000 191.320000 350.100000 ;
        RECT 190.120000 355.060000 191.320000 355.540000 ;
        RECT 190.120000 376.820000 191.320000 377.300000 ;
        RECT 190.120000 371.380000 191.320000 371.860000 ;
        RECT 190.120000 365.940000 191.320000 366.420000 ;
        RECT 145.120000 382.260000 146.320000 382.740000 ;
        RECT 145.120000 387.700000 146.320000 388.180000 ;
        RECT 145.120000 393.140000 146.320000 393.620000 ;
        RECT 145.120000 409.460000 146.320000 409.940000 ;
        RECT 145.120000 404.020000 146.320000 404.500000 ;
        RECT 145.120000 398.580000 146.320000 399.060000 ;
        RECT 190.120000 382.260000 191.320000 382.740000 ;
        RECT 190.120000 387.700000 191.320000 388.180000 ;
        RECT 190.120000 393.140000 191.320000 393.620000 ;
        RECT 190.120000 409.460000 191.320000 409.940000 ;
        RECT 190.120000 404.020000 191.320000 404.500000 ;
        RECT 190.120000 398.580000 191.320000 399.060000 ;
        RECT 235.120000 360.500000 236.320000 360.980000 ;
        RECT 235.120000 355.060000 236.320000 355.540000 ;
        RECT 235.120000 349.620000 236.320000 350.100000 ;
        RECT 235.120000 344.180000 236.320000 344.660000 ;
        RECT 235.120000 376.820000 236.320000 377.300000 ;
        RECT 235.120000 371.380000 236.320000 371.860000 ;
        RECT 235.120000 365.940000 236.320000 366.420000 ;
        RECT 235.120000 393.140000 236.320000 393.620000 ;
        RECT 235.120000 387.700000 236.320000 388.180000 ;
        RECT 235.120000 382.260000 236.320000 382.740000 ;
        RECT 235.120000 409.460000 236.320000 409.940000 ;
        RECT 235.120000 398.580000 236.320000 399.060000 ;
        RECT 235.120000 404.020000 236.320000 404.500000 ;
        RECT 2.560000 420.340000 4.560000 420.820000 ;
        RECT 9.955000 420.340000 11.320000 420.820000 ;
        RECT 2.560000 414.900000 4.560000 415.380000 ;
        RECT 9.955000 414.900000 11.320000 415.380000 ;
        RECT 2.560000 425.780000 4.560000 426.260000 ;
        RECT 9.955000 425.780000 11.320000 426.260000 ;
        RECT 2.560000 436.660000 4.560000 437.140000 ;
        RECT 9.955000 436.660000 11.320000 437.140000 ;
        RECT 2.560000 431.220000 4.560000 431.700000 ;
        RECT 9.955000 431.220000 11.320000 431.700000 ;
        RECT 2.560000 442.100000 4.560000 442.580000 ;
        RECT 9.955000 442.100000 11.320000 442.580000 ;
        RECT 55.120000 414.900000 56.320000 415.380000 ;
        RECT 55.120000 420.340000 56.320000 420.820000 ;
        RECT 55.120000 425.780000 56.320000 426.260000 ;
        RECT 55.120000 442.100000 56.320000 442.580000 ;
        RECT 55.120000 436.660000 56.320000 437.140000 ;
        RECT 55.120000 431.220000 56.320000 431.700000 ;
        RECT 2.560000 463.860000 4.560000 464.340000 ;
        RECT 9.955000 463.860000 11.320000 464.340000 ;
        RECT 2.560000 452.980000 4.560000 453.460000 ;
        RECT 9.955000 452.980000 11.320000 453.460000 ;
        RECT 2.560000 447.540000 4.560000 448.020000 ;
        RECT 9.955000 447.540000 11.320000 448.020000 ;
        RECT 2.560000 458.420000 4.560000 458.900000 ;
        RECT 9.955000 458.420000 11.320000 458.900000 ;
        RECT 2.560000 469.300000 4.560000 469.780000 ;
        RECT 9.955000 469.300000 11.320000 469.780000 ;
        RECT 2.560000 480.180000 4.560000 480.660000 ;
        RECT 9.955000 480.180000 11.320000 480.660000 ;
        RECT 2.560000 474.740000 4.560000 475.220000 ;
        RECT 9.955000 474.740000 11.320000 475.220000 ;
        RECT 55.120000 463.860000 56.320000 464.340000 ;
        RECT 55.120000 447.540000 56.320000 448.020000 ;
        RECT 55.120000 452.980000 56.320000 453.460000 ;
        RECT 55.120000 458.420000 56.320000 458.900000 ;
        RECT 55.120000 480.180000 56.320000 480.660000 ;
        RECT 55.120000 474.740000 56.320000 475.220000 ;
        RECT 55.120000 469.300000 56.320000 469.780000 ;
        RECT 100.120000 442.100000 101.320000 442.580000 ;
        RECT 100.120000 436.660000 101.320000 437.140000 ;
        RECT 100.120000 414.900000 101.320000 415.380000 ;
        RECT 100.120000 420.340000 101.320000 420.820000 ;
        RECT 100.120000 425.780000 101.320000 426.260000 ;
        RECT 100.120000 431.220000 101.320000 431.700000 ;
        RECT 100.120000 480.180000 101.320000 480.660000 ;
        RECT 100.120000 474.740000 101.320000 475.220000 ;
        RECT 100.120000 469.300000 101.320000 469.780000 ;
        RECT 100.120000 447.540000 101.320000 448.020000 ;
        RECT 100.120000 452.980000 101.320000 453.460000 ;
        RECT 100.120000 458.420000 101.320000 458.900000 ;
        RECT 100.120000 463.860000 101.320000 464.340000 ;
        RECT 2.560000 485.620000 4.560000 486.100000 ;
        RECT 9.955000 485.620000 11.320000 486.100000 ;
        RECT 2.560000 496.500000 4.560000 496.980000 ;
        RECT 9.955000 496.500000 11.320000 496.980000 ;
        RECT 2.560000 491.060000 4.560000 491.540000 ;
        RECT 9.955000 491.060000 11.320000 491.540000 ;
        RECT 2.560000 501.940000 4.560000 502.420000 ;
        RECT 9.955000 501.940000 11.320000 502.420000 ;
        RECT 2.560000 512.820000 4.560000 513.300000 ;
        RECT 9.955000 512.820000 11.320000 513.300000 ;
        RECT 2.560000 507.380000 4.560000 507.860000 ;
        RECT 9.955000 507.380000 11.320000 507.860000 ;
        RECT 55.120000 485.620000 56.320000 486.100000 ;
        RECT 55.120000 491.060000 56.320000 491.540000 ;
        RECT 55.120000 496.500000 56.320000 496.980000 ;
        RECT 55.120000 512.820000 56.320000 513.300000 ;
        RECT 55.120000 507.380000 56.320000 507.860000 ;
        RECT 55.120000 501.940000 56.320000 502.420000 ;
        RECT 2.560000 523.700000 4.560000 524.180000 ;
        RECT 9.955000 523.700000 11.320000 524.180000 ;
        RECT 2.560000 518.260000 4.560000 518.740000 ;
        RECT 9.955000 518.260000 11.320000 518.740000 ;
        RECT 2.560000 529.140000 4.560000 529.620000 ;
        RECT 9.955000 529.140000 11.320000 529.620000 ;
        RECT 2.560000 534.580000 4.560000 535.060000 ;
        RECT 9.955000 534.580000 11.320000 535.060000 ;
        RECT 55.120000 534.580000 56.320000 535.060000 ;
        RECT 55.120000 529.140000 56.320000 529.620000 ;
        RECT 55.120000 523.700000 56.320000 524.180000 ;
        RECT 55.120000 518.260000 56.320000 518.740000 ;
        RECT 100.120000 512.820000 101.320000 513.300000 ;
        RECT 100.120000 507.380000 101.320000 507.860000 ;
        RECT 100.120000 485.620000 101.320000 486.100000 ;
        RECT 100.120000 491.060000 101.320000 491.540000 ;
        RECT 100.120000 496.500000 101.320000 496.980000 ;
        RECT 100.120000 501.940000 101.320000 502.420000 ;
        RECT 100.120000 534.580000 101.320000 535.060000 ;
        RECT 100.120000 529.140000 101.320000 529.620000 ;
        RECT 100.120000 523.700000 101.320000 524.180000 ;
        RECT 100.120000 518.260000 101.320000 518.740000 ;
        RECT 145.120000 414.900000 146.320000 415.380000 ;
        RECT 145.120000 420.340000 146.320000 420.820000 ;
        RECT 145.120000 425.780000 146.320000 426.260000 ;
        RECT 145.120000 442.100000 146.320000 442.580000 ;
        RECT 145.120000 436.660000 146.320000 437.140000 ;
        RECT 145.120000 431.220000 146.320000 431.700000 ;
        RECT 190.120000 414.900000 191.320000 415.380000 ;
        RECT 190.120000 420.340000 191.320000 420.820000 ;
        RECT 190.120000 425.780000 191.320000 426.260000 ;
        RECT 190.120000 442.100000 191.320000 442.580000 ;
        RECT 190.120000 436.660000 191.320000 437.140000 ;
        RECT 190.120000 431.220000 191.320000 431.700000 ;
        RECT 145.120000 463.860000 146.320000 464.340000 ;
        RECT 145.120000 447.540000 146.320000 448.020000 ;
        RECT 145.120000 452.980000 146.320000 453.460000 ;
        RECT 145.120000 458.420000 146.320000 458.900000 ;
        RECT 145.120000 480.180000 146.320000 480.660000 ;
        RECT 145.120000 474.740000 146.320000 475.220000 ;
        RECT 145.120000 469.300000 146.320000 469.780000 ;
        RECT 190.120000 463.860000 191.320000 464.340000 ;
        RECT 190.120000 447.540000 191.320000 448.020000 ;
        RECT 190.120000 452.980000 191.320000 453.460000 ;
        RECT 190.120000 458.420000 191.320000 458.900000 ;
        RECT 190.120000 480.180000 191.320000 480.660000 ;
        RECT 190.120000 474.740000 191.320000 475.220000 ;
        RECT 190.120000 469.300000 191.320000 469.780000 ;
        RECT 235.120000 425.780000 236.320000 426.260000 ;
        RECT 235.120000 420.340000 236.320000 420.820000 ;
        RECT 235.120000 414.900000 236.320000 415.380000 ;
        RECT 235.120000 442.100000 236.320000 442.580000 ;
        RECT 235.120000 431.220000 236.320000 431.700000 ;
        RECT 235.120000 436.660000 236.320000 437.140000 ;
        RECT 235.120000 463.860000 236.320000 464.340000 ;
        RECT 235.120000 458.420000 236.320000 458.900000 ;
        RECT 235.120000 452.980000 236.320000 453.460000 ;
        RECT 235.120000 447.540000 236.320000 448.020000 ;
        RECT 235.120000 480.180000 236.320000 480.660000 ;
        RECT 235.120000 474.740000 236.320000 475.220000 ;
        RECT 235.120000 469.300000 236.320000 469.780000 ;
        RECT 145.120000 485.620000 146.320000 486.100000 ;
        RECT 145.120000 491.060000 146.320000 491.540000 ;
        RECT 145.120000 496.500000 146.320000 496.980000 ;
        RECT 145.120000 512.820000 146.320000 513.300000 ;
        RECT 145.120000 507.380000 146.320000 507.860000 ;
        RECT 145.120000 501.940000 146.320000 502.420000 ;
        RECT 190.120000 485.620000 191.320000 486.100000 ;
        RECT 190.120000 491.060000 191.320000 491.540000 ;
        RECT 190.120000 496.500000 191.320000 496.980000 ;
        RECT 190.120000 512.820000 191.320000 513.300000 ;
        RECT 190.120000 507.380000 191.320000 507.860000 ;
        RECT 190.120000 501.940000 191.320000 502.420000 ;
        RECT 145.120000 534.580000 146.320000 535.060000 ;
        RECT 145.120000 529.140000 146.320000 529.620000 ;
        RECT 145.120000 523.700000 146.320000 524.180000 ;
        RECT 145.120000 518.260000 146.320000 518.740000 ;
        RECT 190.120000 534.580000 191.320000 535.060000 ;
        RECT 190.120000 529.140000 191.320000 529.620000 ;
        RECT 190.120000 523.700000 191.320000 524.180000 ;
        RECT 190.120000 518.260000 191.320000 518.740000 ;
        RECT 235.120000 496.500000 236.320000 496.980000 ;
        RECT 235.120000 491.060000 236.320000 491.540000 ;
        RECT 235.120000 485.620000 236.320000 486.100000 ;
        RECT 235.120000 512.820000 236.320000 513.300000 ;
        RECT 235.120000 501.940000 236.320000 502.420000 ;
        RECT 235.120000 507.380000 236.320000 507.860000 ;
        RECT 235.120000 534.580000 236.320000 535.060000 ;
        RECT 235.120000 529.140000 236.320000 529.620000 ;
        RECT 235.120000 523.700000 236.320000 524.180000 ;
        RECT 235.120000 518.260000 236.320000 518.740000 ;
        RECT 280.120000 278.900000 281.320000 279.380000 ;
        RECT 280.120000 284.340000 281.320000 284.820000 ;
        RECT 280.120000 289.780000 281.320000 290.260000 ;
        RECT 280.120000 306.100000 281.320000 306.580000 ;
        RECT 280.120000 300.660000 281.320000 301.140000 ;
        RECT 280.120000 295.220000 281.320000 295.700000 ;
        RECT 325.120000 278.900000 326.320000 279.380000 ;
        RECT 325.120000 284.340000 326.320000 284.820000 ;
        RECT 325.120000 289.780000 326.320000 290.260000 ;
        RECT 325.120000 306.100000 326.320000 306.580000 ;
        RECT 325.120000 300.660000 326.320000 301.140000 ;
        RECT 325.120000 295.220000 326.320000 295.700000 ;
        RECT 280.120000 311.540000 281.320000 312.020000 ;
        RECT 280.120000 316.980000 281.320000 317.460000 ;
        RECT 280.120000 322.420000 281.320000 322.900000 ;
        RECT 280.120000 338.740000 281.320000 339.220000 ;
        RECT 280.120000 333.300000 281.320000 333.780000 ;
        RECT 280.120000 327.860000 281.320000 328.340000 ;
        RECT 325.120000 311.540000 326.320000 312.020000 ;
        RECT 325.120000 316.980000 326.320000 317.460000 ;
        RECT 325.120000 322.420000 326.320000 322.900000 ;
        RECT 325.120000 338.740000 326.320000 339.220000 ;
        RECT 325.120000 333.300000 326.320000 333.780000 ;
        RECT 325.120000 327.860000 326.320000 328.340000 ;
        RECT 370.120000 289.780000 371.320000 290.260000 ;
        RECT 370.120000 284.340000 371.320000 284.820000 ;
        RECT 370.120000 278.900000 371.320000 279.380000 ;
        RECT 370.120000 306.100000 371.320000 306.580000 ;
        RECT 370.120000 295.220000 371.320000 295.700000 ;
        RECT 370.120000 300.660000 371.320000 301.140000 ;
        RECT 370.120000 322.420000 371.320000 322.900000 ;
        RECT 370.120000 316.980000 371.320000 317.460000 ;
        RECT 370.120000 311.540000 371.320000 312.020000 ;
        RECT 370.120000 338.740000 371.320000 339.220000 ;
        RECT 370.120000 327.860000 371.320000 328.340000 ;
        RECT 370.120000 333.300000 371.320000 333.780000 ;
        RECT 280.120000 360.500000 281.320000 360.980000 ;
        RECT 280.120000 344.180000 281.320000 344.660000 ;
        RECT 280.120000 349.620000 281.320000 350.100000 ;
        RECT 280.120000 355.060000 281.320000 355.540000 ;
        RECT 280.120000 376.820000 281.320000 377.300000 ;
        RECT 280.120000 371.380000 281.320000 371.860000 ;
        RECT 280.120000 365.940000 281.320000 366.420000 ;
        RECT 325.120000 360.500000 326.320000 360.980000 ;
        RECT 325.120000 344.180000 326.320000 344.660000 ;
        RECT 325.120000 349.620000 326.320000 350.100000 ;
        RECT 325.120000 355.060000 326.320000 355.540000 ;
        RECT 325.120000 376.820000 326.320000 377.300000 ;
        RECT 325.120000 371.380000 326.320000 371.860000 ;
        RECT 325.120000 365.940000 326.320000 366.420000 ;
        RECT 280.120000 382.260000 281.320000 382.740000 ;
        RECT 280.120000 387.700000 281.320000 388.180000 ;
        RECT 280.120000 393.140000 281.320000 393.620000 ;
        RECT 280.120000 409.460000 281.320000 409.940000 ;
        RECT 280.120000 404.020000 281.320000 404.500000 ;
        RECT 280.120000 398.580000 281.320000 399.060000 ;
        RECT 325.120000 382.260000 326.320000 382.740000 ;
        RECT 325.120000 387.700000 326.320000 388.180000 ;
        RECT 325.120000 393.140000 326.320000 393.620000 ;
        RECT 325.120000 409.460000 326.320000 409.940000 ;
        RECT 325.120000 404.020000 326.320000 404.500000 ;
        RECT 325.120000 398.580000 326.320000 399.060000 ;
        RECT 370.120000 360.500000 371.320000 360.980000 ;
        RECT 370.120000 355.060000 371.320000 355.540000 ;
        RECT 370.120000 349.620000 371.320000 350.100000 ;
        RECT 370.120000 344.180000 371.320000 344.660000 ;
        RECT 370.120000 376.820000 371.320000 377.300000 ;
        RECT 370.120000 371.380000 371.320000 371.860000 ;
        RECT 370.120000 365.940000 371.320000 366.420000 ;
        RECT 370.120000 393.140000 371.320000 393.620000 ;
        RECT 370.120000 387.700000 371.320000 388.180000 ;
        RECT 370.120000 382.260000 371.320000 382.740000 ;
        RECT 370.120000 409.460000 371.320000 409.940000 ;
        RECT 370.120000 398.580000 371.320000 399.060000 ;
        RECT 370.120000 404.020000 371.320000 404.500000 ;
        RECT 415.120000 278.900000 416.320000 279.380000 ;
        RECT 415.120000 284.340000 416.320000 284.820000 ;
        RECT 415.120000 289.780000 416.320000 290.260000 ;
        RECT 415.120000 306.100000 416.320000 306.580000 ;
        RECT 415.120000 300.660000 416.320000 301.140000 ;
        RECT 415.120000 295.220000 416.320000 295.700000 ;
        RECT 460.120000 278.900000 461.320000 279.380000 ;
        RECT 460.120000 284.340000 461.320000 284.820000 ;
        RECT 460.120000 289.780000 461.320000 290.260000 ;
        RECT 460.120000 306.100000 461.320000 306.580000 ;
        RECT 460.120000 300.660000 461.320000 301.140000 ;
        RECT 460.120000 295.220000 461.320000 295.700000 ;
        RECT 415.120000 311.540000 416.320000 312.020000 ;
        RECT 415.120000 316.980000 416.320000 317.460000 ;
        RECT 415.120000 322.420000 416.320000 322.900000 ;
        RECT 415.120000 338.740000 416.320000 339.220000 ;
        RECT 415.120000 333.300000 416.320000 333.780000 ;
        RECT 415.120000 327.860000 416.320000 328.340000 ;
        RECT 460.120000 311.540000 461.320000 312.020000 ;
        RECT 460.120000 316.980000 461.320000 317.460000 ;
        RECT 460.120000 322.420000 461.320000 322.900000 ;
        RECT 460.120000 338.740000 461.320000 339.220000 ;
        RECT 460.120000 333.300000 461.320000 333.780000 ;
        RECT 460.120000 327.860000 461.320000 328.340000 ;
        RECT 505.120000 289.780000 506.320000 290.260000 ;
        RECT 505.120000 284.340000 506.320000 284.820000 ;
        RECT 505.120000 278.900000 506.320000 279.380000 ;
        RECT 505.120000 306.100000 506.320000 306.580000 ;
        RECT 505.120000 295.220000 506.320000 295.700000 ;
        RECT 505.120000 300.660000 506.320000 301.140000 ;
        RECT 545.600000 289.780000 547.600000 290.260000 ;
        RECT 545.600000 278.900000 547.600000 279.380000 ;
        RECT 545.600000 284.340000 547.600000 284.820000 ;
        RECT 545.600000 306.100000 547.600000 306.580000 ;
        RECT 545.600000 300.660000 547.600000 301.140000 ;
        RECT 545.600000 295.220000 547.600000 295.700000 ;
        RECT 505.120000 322.420000 506.320000 322.900000 ;
        RECT 505.120000 316.980000 506.320000 317.460000 ;
        RECT 505.120000 311.540000 506.320000 312.020000 ;
        RECT 505.120000 338.740000 506.320000 339.220000 ;
        RECT 505.120000 327.860000 506.320000 328.340000 ;
        RECT 505.120000 333.300000 506.320000 333.780000 ;
        RECT 545.600000 322.420000 547.600000 322.900000 ;
        RECT 545.600000 311.540000 547.600000 312.020000 ;
        RECT 545.600000 316.980000 547.600000 317.460000 ;
        RECT 545.600000 338.740000 547.600000 339.220000 ;
        RECT 545.600000 333.300000 547.600000 333.780000 ;
        RECT 545.600000 327.860000 547.600000 328.340000 ;
        RECT 415.120000 360.500000 416.320000 360.980000 ;
        RECT 415.120000 344.180000 416.320000 344.660000 ;
        RECT 415.120000 349.620000 416.320000 350.100000 ;
        RECT 415.120000 355.060000 416.320000 355.540000 ;
        RECT 415.120000 376.820000 416.320000 377.300000 ;
        RECT 415.120000 371.380000 416.320000 371.860000 ;
        RECT 415.120000 365.940000 416.320000 366.420000 ;
        RECT 460.120000 360.500000 461.320000 360.980000 ;
        RECT 460.120000 344.180000 461.320000 344.660000 ;
        RECT 460.120000 349.620000 461.320000 350.100000 ;
        RECT 460.120000 355.060000 461.320000 355.540000 ;
        RECT 460.120000 376.820000 461.320000 377.300000 ;
        RECT 460.120000 371.380000 461.320000 371.860000 ;
        RECT 460.120000 365.940000 461.320000 366.420000 ;
        RECT 415.120000 382.260000 416.320000 382.740000 ;
        RECT 415.120000 387.700000 416.320000 388.180000 ;
        RECT 415.120000 393.140000 416.320000 393.620000 ;
        RECT 415.120000 409.460000 416.320000 409.940000 ;
        RECT 415.120000 404.020000 416.320000 404.500000 ;
        RECT 415.120000 398.580000 416.320000 399.060000 ;
        RECT 460.120000 382.260000 461.320000 382.740000 ;
        RECT 460.120000 387.700000 461.320000 388.180000 ;
        RECT 460.120000 393.140000 461.320000 393.620000 ;
        RECT 460.120000 409.460000 461.320000 409.940000 ;
        RECT 460.120000 404.020000 461.320000 404.500000 ;
        RECT 460.120000 398.580000 461.320000 399.060000 ;
        RECT 505.120000 360.500000 506.320000 360.980000 ;
        RECT 505.120000 355.060000 506.320000 355.540000 ;
        RECT 505.120000 349.620000 506.320000 350.100000 ;
        RECT 505.120000 344.180000 506.320000 344.660000 ;
        RECT 505.120000 376.820000 506.320000 377.300000 ;
        RECT 505.120000 371.380000 506.320000 371.860000 ;
        RECT 505.120000 365.940000 506.320000 366.420000 ;
        RECT 545.600000 360.500000 547.600000 360.980000 ;
        RECT 545.600000 355.060000 547.600000 355.540000 ;
        RECT 545.600000 344.180000 547.600000 344.660000 ;
        RECT 545.600000 349.620000 547.600000 350.100000 ;
        RECT 545.600000 376.820000 547.600000 377.300000 ;
        RECT 545.600000 371.380000 547.600000 371.860000 ;
        RECT 545.600000 365.940000 547.600000 366.420000 ;
        RECT 505.120000 393.140000 506.320000 393.620000 ;
        RECT 505.120000 387.700000 506.320000 388.180000 ;
        RECT 505.120000 382.260000 506.320000 382.740000 ;
        RECT 505.120000 409.460000 506.320000 409.940000 ;
        RECT 505.120000 398.580000 506.320000 399.060000 ;
        RECT 505.120000 404.020000 506.320000 404.500000 ;
        RECT 545.600000 393.140000 547.600000 393.620000 ;
        RECT 545.600000 382.260000 547.600000 382.740000 ;
        RECT 545.600000 387.700000 547.600000 388.180000 ;
        RECT 545.600000 409.460000 547.600000 409.940000 ;
        RECT 545.600000 404.020000 547.600000 404.500000 ;
        RECT 545.600000 398.580000 547.600000 399.060000 ;
        RECT 280.120000 414.900000 281.320000 415.380000 ;
        RECT 280.120000 420.340000 281.320000 420.820000 ;
        RECT 280.120000 425.780000 281.320000 426.260000 ;
        RECT 280.120000 442.100000 281.320000 442.580000 ;
        RECT 280.120000 436.660000 281.320000 437.140000 ;
        RECT 280.120000 431.220000 281.320000 431.700000 ;
        RECT 325.120000 414.900000 326.320000 415.380000 ;
        RECT 325.120000 420.340000 326.320000 420.820000 ;
        RECT 325.120000 425.780000 326.320000 426.260000 ;
        RECT 325.120000 442.100000 326.320000 442.580000 ;
        RECT 325.120000 436.660000 326.320000 437.140000 ;
        RECT 325.120000 431.220000 326.320000 431.700000 ;
        RECT 280.120000 463.860000 281.320000 464.340000 ;
        RECT 280.120000 447.540000 281.320000 448.020000 ;
        RECT 280.120000 452.980000 281.320000 453.460000 ;
        RECT 280.120000 458.420000 281.320000 458.900000 ;
        RECT 280.120000 480.180000 281.320000 480.660000 ;
        RECT 280.120000 474.740000 281.320000 475.220000 ;
        RECT 280.120000 469.300000 281.320000 469.780000 ;
        RECT 325.120000 463.860000 326.320000 464.340000 ;
        RECT 325.120000 447.540000 326.320000 448.020000 ;
        RECT 325.120000 452.980000 326.320000 453.460000 ;
        RECT 325.120000 458.420000 326.320000 458.900000 ;
        RECT 325.120000 480.180000 326.320000 480.660000 ;
        RECT 325.120000 474.740000 326.320000 475.220000 ;
        RECT 325.120000 469.300000 326.320000 469.780000 ;
        RECT 370.120000 425.780000 371.320000 426.260000 ;
        RECT 370.120000 420.340000 371.320000 420.820000 ;
        RECT 370.120000 414.900000 371.320000 415.380000 ;
        RECT 370.120000 442.100000 371.320000 442.580000 ;
        RECT 370.120000 431.220000 371.320000 431.700000 ;
        RECT 370.120000 436.660000 371.320000 437.140000 ;
        RECT 370.120000 463.860000 371.320000 464.340000 ;
        RECT 370.120000 458.420000 371.320000 458.900000 ;
        RECT 370.120000 452.980000 371.320000 453.460000 ;
        RECT 370.120000 447.540000 371.320000 448.020000 ;
        RECT 370.120000 480.180000 371.320000 480.660000 ;
        RECT 370.120000 474.740000 371.320000 475.220000 ;
        RECT 370.120000 469.300000 371.320000 469.780000 ;
        RECT 280.120000 485.620000 281.320000 486.100000 ;
        RECT 280.120000 491.060000 281.320000 491.540000 ;
        RECT 280.120000 496.500000 281.320000 496.980000 ;
        RECT 280.120000 512.820000 281.320000 513.300000 ;
        RECT 280.120000 507.380000 281.320000 507.860000 ;
        RECT 280.120000 501.940000 281.320000 502.420000 ;
        RECT 325.120000 485.620000 326.320000 486.100000 ;
        RECT 325.120000 491.060000 326.320000 491.540000 ;
        RECT 325.120000 496.500000 326.320000 496.980000 ;
        RECT 325.120000 512.820000 326.320000 513.300000 ;
        RECT 325.120000 507.380000 326.320000 507.860000 ;
        RECT 325.120000 501.940000 326.320000 502.420000 ;
        RECT 280.120000 534.580000 281.320000 535.060000 ;
        RECT 280.120000 529.140000 281.320000 529.620000 ;
        RECT 280.120000 523.700000 281.320000 524.180000 ;
        RECT 280.120000 518.260000 281.320000 518.740000 ;
        RECT 325.120000 534.580000 326.320000 535.060000 ;
        RECT 325.120000 529.140000 326.320000 529.620000 ;
        RECT 325.120000 523.700000 326.320000 524.180000 ;
        RECT 325.120000 518.260000 326.320000 518.740000 ;
        RECT 370.120000 496.500000 371.320000 496.980000 ;
        RECT 370.120000 491.060000 371.320000 491.540000 ;
        RECT 370.120000 485.620000 371.320000 486.100000 ;
        RECT 370.120000 512.820000 371.320000 513.300000 ;
        RECT 370.120000 501.940000 371.320000 502.420000 ;
        RECT 370.120000 507.380000 371.320000 507.860000 ;
        RECT 370.120000 534.580000 371.320000 535.060000 ;
        RECT 370.120000 529.140000 371.320000 529.620000 ;
        RECT 370.120000 523.700000 371.320000 524.180000 ;
        RECT 370.120000 518.260000 371.320000 518.740000 ;
        RECT 415.120000 414.900000 416.320000 415.380000 ;
        RECT 415.120000 420.340000 416.320000 420.820000 ;
        RECT 415.120000 425.780000 416.320000 426.260000 ;
        RECT 415.120000 442.100000 416.320000 442.580000 ;
        RECT 415.120000 436.660000 416.320000 437.140000 ;
        RECT 415.120000 431.220000 416.320000 431.700000 ;
        RECT 460.120000 414.900000 461.320000 415.380000 ;
        RECT 460.120000 420.340000 461.320000 420.820000 ;
        RECT 460.120000 425.780000 461.320000 426.260000 ;
        RECT 460.120000 442.100000 461.320000 442.580000 ;
        RECT 460.120000 436.660000 461.320000 437.140000 ;
        RECT 460.120000 431.220000 461.320000 431.700000 ;
        RECT 415.120000 463.860000 416.320000 464.340000 ;
        RECT 415.120000 447.540000 416.320000 448.020000 ;
        RECT 415.120000 452.980000 416.320000 453.460000 ;
        RECT 415.120000 458.420000 416.320000 458.900000 ;
        RECT 415.120000 480.180000 416.320000 480.660000 ;
        RECT 415.120000 474.740000 416.320000 475.220000 ;
        RECT 415.120000 469.300000 416.320000 469.780000 ;
        RECT 460.120000 463.860000 461.320000 464.340000 ;
        RECT 460.120000 447.540000 461.320000 448.020000 ;
        RECT 460.120000 452.980000 461.320000 453.460000 ;
        RECT 460.120000 458.420000 461.320000 458.900000 ;
        RECT 460.120000 480.180000 461.320000 480.660000 ;
        RECT 460.120000 474.740000 461.320000 475.220000 ;
        RECT 460.120000 469.300000 461.320000 469.780000 ;
        RECT 505.120000 425.780000 506.320000 426.260000 ;
        RECT 505.120000 420.340000 506.320000 420.820000 ;
        RECT 505.120000 414.900000 506.320000 415.380000 ;
        RECT 505.120000 442.100000 506.320000 442.580000 ;
        RECT 505.120000 431.220000 506.320000 431.700000 ;
        RECT 505.120000 436.660000 506.320000 437.140000 ;
        RECT 545.600000 425.780000 547.600000 426.260000 ;
        RECT 545.600000 414.900000 547.600000 415.380000 ;
        RECT 545.600000 420.340000 547.600000 420.820000 ;
        RECT 545.600000 442.100000 547.600000 442.580000 ;
        RECT 545.600000 436.660000 547.600000 437.140000 ;
        RECT 545.600000 431.220000 547.600000 431.700000 ;
        RECT 505.120000 463.860000 506.320000 464.340000 ;
        RECT 505.120000 458.420000 506.320000 458.900000 ;
        RECT 505.120000 452.980000 506.320000 453.460000 ;
        RECT 505.120000 447.540000 506.320000 448.020000 ;
        RECT 505.120000 480.180000 506.320000 480.660000 ;
        RECT 505.120000 474.740000 506.320000 475.220000 ;
        RECT 505.120000 469.300000 506.320000 469.780000 ;
        RECT 545.600000 463.860000 547.600000 464.340000 ;
        RECT 545.600000 458.420000 547.600000 458.900000 ;
        RECT 545.600000 447.540000 547.600000 448.020000 ;
        RECT 545.600000 452.980000 547.600000 453.460000 ;
        RECT 545.600000 480.180000 547.600000 480.660000 ;
        RECT 545.600000 474.740000 547.600000 475.220000 ;
        RECT 545.600000 469.300000 547.600000 469.780000 ;
        RECT 415.120000 485.620000 416.320000 486.100000 ;
        RECT 415.120000 491.060000 416.320000 491.540000 ;
        RECT 415.120000 496.500000 416.320000 496.980000 ;
        RECT 415.120000 512.820000 416.320000 513.300000 ;
        RECT 415.120000 507.380000 416.320000 507.860000 ;
        RECT 415.120000 501.940000 416.320000 502.420000 ;
        RECT 460.120000 485.620000 461.320000 486.100000 ;
        RECT 460.120000 491.060000 461.320000 491.540000 ;
        RECT 460.120000 496.500000 461.320000 496.980000 ;
        RECT 460.120000 512.820000 461.320000 513.300000 ;
        RECT 460.120000 507.380000 461.320000 507.860000 ;
        RECT 460.120000 501.940000 461.320000 502.420000 ;
        RECT 415.120000 534.580000 416.320000 535.060000 ;
        RECT 415.120000 529.140000 416.320000 529.620000 ;
        RECT 415.120000 523.700000 416.320000 524.180000 ;
        RECT 415.120000 518.260000 416.320000 518.740000 ;
        RECT 460.120000 534.580000 461.320000 535.060000 ;
        RECT 460.120000 529.140000 461.320000 529.620000 ;
        RECT 460.120000 523.700000 461.320000 524.180000 ;
        RECT 460.120000 518.260000 461.320000 518.740000 ;
        RECT 505.120000 496.500000 506.320000 496.980000 ;
        RECT 505.120000 491.060000 506.320000 491.540000 ;
        RECT 505.120000 485.620000 506.320000 486.100000 ;
        RECT 505.120000 512.820000 506.320000 513.300000 ;
        RECT 505.120000 501.940000 506.320000 502.420000 ;
        RECT 505.120000 507.380000 506.320000 507.860000 ;
        RECT 545.600000 496.500000 547.600000 496.980000 ;
        RECT 545.600000 485.620000 547.600000 486.100000 ;
        RECT 545.600000 491.060000 547.600000 491.540000 ;
        RECT 545.600000 512.820000 547.600000 513.300000 ;
        RECT 545.600000 507.380000 547.600000 507.860000 ;
        RECT 545.600000 501.940000 547.600000 502.420000 ;
        RECT 505.120000 518.260000 506.320000 518.740000 ;
        RECT 505.120000 523.700000 506.320000 524.180000 ;
        RECT 505.120000 529.140000 506.320000 529.620000 ;
        RECT 505.120000 534.580000 506.320000 535.060000 ;
        RECT 545.600000 518.260000 547.600000 518.740000 ;
        RECT 545.600000 523.700000 547.600000 524.180000 ;
        RECT 545.600000 529.140000 547.600000 529.620000 ;
        RECT 545.600000 534.580000 547.600000 535.060000 ;
      LAYER met4 ;
        RECT 505.120000 2.430000 506.320000 546.160000 ;
        RECT 460.120000 2.430000 461.320000 546.160000 ;
        RECT 415.120000 2.430000 416.320000 546.160000 ;
        RECT 370.120000 2.430000 371.320000 546.160000 ;
        RECT 325.120000 2.430000 326.320000 546.160000 ;
        RECT 280.120000 2.430000 281.320000 546.160000 ;
        RECT 235.120000 2.430000 236.320000 546.160000 ;
        RECT 190.120000 2.430000 191.320000 546.160000 ;
        RECT 145.120000 2.430000 146.320000 546.160000 ;
        RECT 100.120000 2.430000 101.320000 546.160000 ;
        RECT 55.120000 2.430000 56.320000 546.160000 ;
        RECT 10.120000 2.430000 11.320000 546.160000 ;
        RECT 545.600000 0.000000 547.600000 549.780000 ;
        RECT 2.560000 0.000000 4.560000 549.780000 ;
        RECT 9.955000 34.100000 11.320000 34.580000 ;
        RECT 9.955000 12.340000 11.320000 12.820000 ;
        RECT 9.955000 23.220000 11.320000 23.700000 ;
        RECT 9.955000 17.780000 11.320000 18.260000 ;
        RECT 9.955000 28.660000 11.320000 29.140000 ;
        RECT 9.955000 39.540000 11.320000 40.020000 ;
        RECT 9.955000 50.420000 11.320000 50.900000 ;
        RECT 9.955000 44.980000 11.320000 45.460000 ;
        RECT 9.955000 55.860000 11.320000 56.340000 ;
        RECT 9.955000 66.740000 11.320000 67.220000 ;
        RECT 9.955000 61.300000 11.320000 61.780000 ;
        RECT 9.955000 72.180000 11.320000 72.660000 ;
        RECT 9.955000 83.060000 11.320000 83.540000 ;
        RECT 9.955000 77.620000 11.320000 78.100000 ;
        RECT 9.955000 93.940000 11.320000 94.420000 ;
        RECT 9.955000 88.500000 11.320000 88.980000 ;
        RECT 9.955000 99.380000 11.320000 99.860000 ;
        RECT 9.955000 110.260000 11.320000 110.740000 ;
        RECT 9.955000 104.820000 11.320000 105.300000 ;
        RECT 9.955000 115.700000 11.320000 116.180000 ;
        RECT 9.955000 126.580000 11.320000 127.060000 ;
        RECT 9.955000 121.140000 11.320000 121.620000 ;
        RECT 9.955000 132.020000 11.320000 132.500000 ;
        RECT 9.955000 142.900000 11.320000 143.380000 ;
        RECT 9.955000 137.460000 11.320000 137.940000 ;
        RECT 9.955000 153.780000 11.320000 154.260000 ;
        RECT 9.955000 148.340000 11.320000 148.820000 ;
        RECT 9.955000 159.220000 11.320000 159.700000 ;
        RECT 9.955000 170.100000 11.320000 170.580000 ;
        RECT 9.955000 164.660000 11.320000 165.140000 ;
        RECT 9.955000 175.540000 11.320000 176.020000 ;
        RECT 9.955000 186.420000 11.320000 186.900000 ;
        RECT 9.955000 180.980000 11.320000 181.460000 ;
        RECT 9.955000 197.300000 11.320000 197.780000 ;
        RECT 9.955000 191.860000 11.320000 192.340000 ;
        RECT 9.955000 202.740000 11.320000 203.220000 ;
        RECT 9.955000 213.620000 11.320000 214.100000 ;
        RECT 9.955000 208.180000 11.320000 208.660000 ;
        RECT 9.955000 219.060000 11.320000 219.540000 ;
        RECT 9.955000 229.940000 11.320000 230.420000 ;
        RECT 9.955000 224.500000 11.320000 224.980000 ;
        RECT 9.955000 235.380000 11.320000 235.860000 ;
        RECT 9.955000 246.260000 11.320000 246.740000 ;
        RECT 9.955000 240.820000 11.320000 241.300000 ;
        RECT 9.955000 257.140000 11.320000 257.620000 ;
        RECT 9.955000 251.700000 11.320000 252.180000 ;
        RECT 9.955000 262.580000 11.320000 263.060000 ;
        RECT 9.955000 273.460000 11.320000 273.940000 ;
        RECT 9.955000 268.020000 11.320000 268.500000 ;
        RECT 9.955000 278.900000 11.320000 279.380000 ;
        RECT 9.955000 289.780000 11.320000 290.260000 ;
        RECT 9.955000 284.340000 11.320000 284.820000 ;
        RECT 9.955000 300.660000 11.320000 301.140000 ;
        RECT 9.955000 295.220000 11.320000 295.700000 ;
        RECT 9.955000 306.100000 11.320000 306.580000 ;
        RECT 9.955000 316.980000 11.320000 317.460000 ;
        RECT 9.955000 311.540000 11.320000 312.020000 ;
        RECT 9.955000 322.420000 11.320000 322.900000 ;
        RECT 9.955000 333.300000 11.320000 333.780000 ;
        RECT 9.955000 327.860000 11.320000 328.340000 ;
        RECT 9.955000 338.740000 11.320000 339.220000 ;
        RECT 9.955000 360.500000 11.320000 360.980000 ;
        RECT 9.955000 349.620000 11.320000 350.100000 ;
        RECT 9.955000 344.180000 11.320000 344.660000 ;
        RECT 9.955000 355.060000 11.320000 355.540000 ;
        RECT 9.955000 365.940000 11.320000 366.420000 ;
        RECT 9.955000 376.820000 11.320000 377.300000 ;
        RECT 9.955000 371.380000 11.320000 371.860000 ;
        RECT 9.955000 382.260000 11.320000 382.740000 ;
        RECT 9.955000 393.140000 11.320000 393.620000 ;
        RECT 9.955000 387.700000 11.320000 388.180000 ;
        RECT 9.955000 398.580000 11.320000 399.060000 ;
        RECT 9.955000 409.460000 11.320000 409.940000 ;
        RECT 9.955000 404.020000 11.320000 404.500000 ;
        RECT 9.955000 420.340000 11.320000 420.820000 ;
        RECT 9.955000 414.900000 11.320000 415.380000 ;
        RECT 9.955000 425.780000 11.320000 426.260000 ;
        RECT 9.955000 436.660000 11.320000 437.140000 ;
        RECT 9.955000 431.220000 11.320000 431.700000 ;
        RECT 9.955000 442.100000 11.320000 442.580000 ;
        RECT 9.955000 463.860000 11.320000 464.340000 ;
        RECT 9.955000 452.980000 11.320000 453.460000 ;
        RECT 9.955000 447.540000 11.320000 448.020000 ;
        RECT 9.955000 458.420000 11.320000 458.900000 ;
        RECT 9.955000 469.300000 11.320000 469.780000 ;
        RECT 9.955000 480.180000 11.320000 480.660000 ;
        RECT 9.955000 474.740000 11.320000 475.220000 ;
        RECT 9.955000 485.620000 11.320000 486.100000 ;
        RECT 9.955000 496.500000 11.320000 496.980000 ;
        RECT 9.955000 491.060000 11.320000 491.540000 ;
        RECT 9.955000 501.940000 11.320000 502.420000 ;
        RECT 9.955000 512.820000 11.320000 513.300000 ;
        RECT 9.955000 507.380000 11.320000 507.860000 ;
        RECT 9.955000 523.700000 11.320000 524.180000 ;
        RECT 9.955000 518.260000 11.320000 518.740000 ;
        RECT 9.955000 529.140000 11.320000 529.620000 ;
        RECT 9.955000 534.580000 11.320000 535.060000 ;
    END
# end of P/G power stripe data as pin

  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 550.160000 549.780000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 550.160000 549.780000 ;
    LAYER met2 ;
      RECT 0.000000 1.040000 550.160000 549.780000 ;
      RECT 539.680000 0.000000 550.160000 1.040000 ;
      RECT 536.920000 0.000000 539.020000 1.040000 ;
      RECT 533.700000 0.000000 536.260000 1.040000 ;
      RECT 530.480000 0.000000 533.040000 1.040000 ;
      RECT 527.260000 0.000000 529.820000 1.040000 ;
      RECT 524.040000 0.000000 526.600000 1.040000 ;
      RECT 520.820000 0.000000 523.380000 1.040000 ;
      RECT 518.060000 0.000000 520.160000 1.040000 ;
      RECT 514.840000 0.000000 517.400000 1.040000 ;
      RECT 511.620000 0.000000 514.180000 1.040000 ;
      RECT 508.400000 0.000000 510.960000 1.040000 ;
      RECT 505.180000 0.000000 507.740000 1.040000 ;
      RECT 501.960000 0.000000 504.520000 1.040000 ;
      RECT 498.740000 0.000000 501.300000 1.040000 ;
      RECT 495.980000 0.000000 498.080000 1.040000 ;
      RECT 492.760000 0.000000 495.320000 1.040000 ;
      RECT 489.540000 0.000000 492.100000 1.040000 ;
      RECT 486.320000 0.000000 488.880000 1.040000 ;
      RECT 483.100000 0.000000 485.660000 1.040000 ;
      RECT 479.880000 0.000000 482.440000 1.040000 ;
      RECT 476.660000 0.000000 479.220000 1.040000 ;
      RECT 473.900000 0.000000 476.000000 1.040000 ;
      RECT 470.680000 0.000000 473.240000 1.040000 ;
      RECT 467.460000 0.000000 470.020000 1.040000 ;
      RECT 464.240000 0.000000 466.800000 1.040000 ;
      RECT 461.020000 0.000000 463.580000 1.040000 ;
      RECT 457.800000 0.000000 460.360000 1.040000 ;
      RECT 455.040000 0.000000 457.140000 1.040000 ;
      RECT 451.820000 0.000000 454.380000 1.040000 ;
      RECT 448.600000 0.000000 451.160000 1.040000 ;
      RECT 445.380000 0.000000 447.940000 1.040000 ;
      RECT 442.160000 0.000000 444.720000 1.040000 ;
      RECT 438.940000 0.000000 441.500000 1.040000 ;
      RECT 435.720000 0.000000 438.280000 1.040000 ;
      RECT 432.960000 0.000000 435.060000 1.040000 ;
      RECT 429.740000 0.000000 432.300000 1.040000 ;
      RECT 426.520000 0.000000 429.080000 1.040000 ;
      RECT 423.300000 0.000000 425.860000 1.040000 ;
      RECT 420.080000 0.000000 422.640000 1.040000 ;
      RECT 416.860000 0.000000 419.420000 1.040000 ;
      RECT 413.640000 0.000000 416.200000 1.040000 ;
      RECT 410.880000 0.000000 412.980000 1.040000 ;
      RECT 407.660000 0.000000 410.220000 1.040000 ;
      RECT 404.440000 0.000000 407.000000 1.040000 ;
      RECT 401.220000 0.000000 403.780000 1.040000 ;
      RECT 398.000000 0.000000 400.560000 1.040000 ;
      RECT 394.780000 0.000000 397.340000 1.040000 ;
      RECT 391.560000 0.000000 394.120000 1.040000 ;
      RECT 388.800000 0.000000 390.900000 1.040000 ;
      RECT 385.580000 0.000000 388.140000 1.040000 ;
      RECT 382.360000 0.000000 384.920000 1.040000 ;
      RECT 379.140000 0.000000 381.700000 1.040000 ;
      RECT 375.920000 0.000000 378.480000 1.040000 ;
      RECT 372.700000 0.000000 375.260000 1.040000 ;
      RECT 369.940000 0.000000 372.040000 1.040000 ;
      RECT 366.720000 0.000000 369.280000 1.040000 ;
      RECT 363.500000 0.000000 366.060000 1.040000 ;
      RECT 360.280000 0.000000 362.840000 1.040000 ;
      RECT 357.060000 0.000000 359.620000 1.040000 ;
      RECT 353.840000 0.000000 356.400000 1.040000 ;
      RECT 350.620000 0.000000 353.180000 1.040000 ;
      RECT 347.860000 0.000000 349.960000 1.040000 ;
      RECT 344.640000 0.000000 347.200000 1.040000 ;
      RECT 341.420000 0.000000 343.980000 1.040000 ;
      RECT 338.200000 0.000000 340.760000 1.040000 ;
      RECT 334.980000 0.000000 337.540000 1.040000 ;
      RECT 331.760000 0.000000 334.320000 1.040000 ;
      RECT 328.540000 0.000000 331.100000 1.040000 ;
      RECT 325.780000 0.000000 327.880000 1.040000 ;
      RECT 322.560000 0.000000 325.120000 1.040000 ;
      RECT 319.340000 0.000000 321.900000 1.040000 ;
      RECT 316.120000 0.000000 318.680000 1.040000 ;
      RECT 312.900000 0.000000 315.460000 1.040000 ;
      RECT 309.680000 0.000000 312.240000 1.040000 ;
      RECT 306.920000 0.000000 309.020000 1.040000 ;
      RECT 303.700000 0.000000 306.260000 1.040000 ;
      RECT 300.480000 0.000000 303.040000 1.040000 ;
      RECT 297.260000 0.000000 299.820000 1.040000 ;
      RECT 294.040000 0.000000 296.600000 1.040000 ;
      RECT 290.820000 0.000000 293.380000 1.040000 ;
      RECT 287.600000 0.000000 290.160000 1.040000 ;
      RECT 284.840000 0.000000 286.940000 1.040000 ;
      RECT 281.620000 0.000000 284.180000 1.040000 ;
      RECT 278.400000 0.000000 280.960000 1.040000 ;
      RECT 275.180000 0.000000 277.740000 1.040000 ;
      RECT 271.960000 0.000000 274.520000 1.040000 ;
      RECT 268.740000 0.000000 271.300000 1.040000 ;
      RECT 265.520000 0.000000 268.080000 1.040000 ;
      RECT 262.760000 0.000000 264.860000 1.040000 ;
      RECT 259.540000 0.000000 262.100000 1.040000 ;
      RECT 256.320000 0.000000 258.880000 1.040000 ;
      RECT 253.100000 0.000000 255.660000 1.040000 ;
      RECT 249.880000 0.000000 252.440000 1.040000 ;
      RECT 246.660000 0.000000 249.220000 1.040000 ;
      RECT 243.440000 0.000000 246.000000 1.040000 ;
      RECT 240.680000 0.000000 242.780000 1.040000 ;
      RECT 237.460000 0.000000 240.020000 1.040000 ;
      RECT 234.240000 0.000000 236.800000 1.040000 ;
      RECT 231.020000 0.000000 233.580000 1.040000 ;
      RECT 227.800000 0.000000 230.360000 1.040000 ;
      RECT 224.580000 0.000000 227.140000 1.040000 ;
      RECT 221.820000 0.000000 223.920000 1.040000 ;
      RECT 218.600000 0.000000 221.160000 1.040000 ;
      RECT 215.380000 0.000000 217.940000 1.040000 ;
      RECT 212.160000 0.000000 214.720000 1.040000 ;
      RECT 208.940000 0.000000 211.500000 1.040000 ;
      RECT 205.720000 0.000000 208.280000 1.040000 ;
      RECT 202.500000 0.000000 205.060000 1.040000 ;
      RECT 199.740000 0.000000 201.840000 1.040000 ;
      RECT 196.520000 0.000000 199.080000 1.040000 ;
      RECT 193.300000 0.000000 195.860000 1.040000 ;
      RECT 190.080000 0.000000 192.640000 1.040000 ;
      RECT 186.860000 0.000000 189.420000 1.040000 ;
      RECT 183.640000 0.000000 186.200000 1.040000 ;
      RECT 180.420000 0.000000 182.980000 1.040000 ;
      RECT 177.660000 0.000000 179.760000 1.040000 ;
      RECT 174.440000 0.000000 177.000000 1.040000 ;
      RECT 171.220000 0.000000 173.780000 1.040000 ;
      RECT 168.000000 0.000000 170.560000 1.040000 ;
      RECT 164.780000 0.000000 167.340000 1.040000 ;
      RECT 161.560000 0.000000 164.120000 1.040000 ;
      RECT 158.800000 0.000000 160.900000 1.040000 ;
      RECT 155.580000 0.000000 158.140000 1.040000 ;
      RECT 152.360000 0.000000 154.920000 1.040000 ;
      RECT 149.140000 0.000000 151.700000 1.040000 ;
      RECT 145.920000 0.000000 148.480000 1.040000 ;
      RECT 142.700000 0.000000 145.260000 1.040000 ;
      RECT 139.480000 0.000000 142.040000 1.040000 ;
      RECT 136.720000 0.000000 138.820000 1.040000 ;
      RECT 133.500000 0.000000 136.060000 1.040000 ;
      RECT 130.280000 0.000000 132.840000 1.040000 ;
      RECT 127.060000 0.000000 129.620000 1.040000 ;
      RECT 123.840000 0.000000 126.400000 1.040000 ;
      RECT 120.620000 0.000000 123.180000 1.040000 ;
      RECT 117.400000 0.000000 119.960000 1.040000 ;
      RECT 114.640000 0.000000 116.740000 1.040000 ;
      RECT 111.420000 0.000000 113.980000 1.040000 ;
      RECT 108.200000 0.000000 110.760000 1.040000 ;
      RECT 104.980000 0.000000 107.540000 1.040000 ;
      RECT 101.760000 0.000000 104.320000 1.040000 ;
      RECT 98.540000 0.000000 101.100000 1.040000 ;
      RECT 95.320000 0.000000 97.880000 1.040000 ;
      RECT 92.560000 0.000000 94.660000 1.040000 ;
      RECT 89.340000 0.000000 91.900000 1.040000 ;
      RECT 86.120000 0.000000 88.680000 1.040000 ;
      RECT 82.900000 0.000000 85.460000 1.040000 ;
      RECT 79.680000 0.000000 82.240000 1.040000 ;
      RECT 76.460000 0.000000 79.020000 1.040000 ;
      RECT 73.700000 0.000000 75.800000 1.040000 ;
      RECT 70.480000 0.000000 73.040000 1.040000 ;
      RECT 67.260000 0.000000 69.820000 1.040000 ;
      RECT 64.040000 0.000000 66.600000 1.040000 ;
      RECT 60.820000 0.000000 63.380000 1.040000 ;
      RECT 57.600000 0.000000 60.160000 1.040000 ;
      RECT 54.380000 0.000000 56.940000 1.040000 ;
      RECT 51.620000 0.000000 53.720000 1.040000 ;
      RECT 48.400000 0.000000 50.960000 1.040000 ;
      RECT 45.180000 0.000000 47.740000 1.040000 ;
      RECT 41.960000 0.000000 44.520000 1.040000 ;
      RECT 38.740000 0.000000 41.300000 1.040000 ;
      RECT 35.520000 0.000000 38.080000 1.040000 ;
      RECT 32.300000 0.000000 34.860000 1.040000 ;
      RECT 29.540000 0.000000 31.640000 1.040000 ;
      RECT 26.320000 0.000000 28.880000 1.040000 ;
      RECT 23.100000 0.000000 25.660000 1.040000 ;
      RECT 19.880000 0.000000 22.440000 1.040000 ;
      RECT 16.660000 0.000000 19.220000 1.040000 ;
      RECT 13.440000 0.000000 16.000000 1.040000 ;
      RECT 10.680000 0.000000 12.780000 1.040000 ;
      RECT 0.000000 0.000000 10.020000 1.040000 ;
    LAYER met3 ;
      RECT 0.000000 546.460000 550.160000 549.780000 ;
      RECT 0.000000 543.460000 550.160000 543.860000 ;
      RECT 0.000000 539.390000 550.160000 540.860000 ;
      RECT 0.000000 538.410000 548.960000 539.390000 ;
      RECT 0.000000 538.080000 550.160000 538.410000 ;
      RECT 544.900000 537.560000 550.160000 538.080000 ;
      RECT 544.900000 537.000000 548.960000 537.560000 ;
      RECT 508.620000 537.000000 542.300000 538.080000 ;
      RECT 463.620000 537.000000 506.820000 538.080000 ;
      RECT 418.620000 537.000000 461.820000 538.080000 ;
      RECT 373.620000 537.000000 416.820000 538.080000 ;
      RECT 328.620000 537.000000 371.820000 538.080000 ;
      RECT 283.620000 537.000000 326.820000 538.080000 ;
      RECT 238.620000 537.000000 281.820000 538.080000 ;
      RECT 193.620000 537.000000 236.820000 538.080000 ;
      RECT 148.620000 537.000000 191.820000 538.080000 ;
      RECT 103.620000 537.000000 146.820000 538.080000 ;
      RECT 58.620000 537.000000 101.820000 538.080000 ;
      RECT 13.620000 537.000000 56.820000 538.080000 ;
      RECT 7.860000 537.000000 11.820000 538.080000 ;
      RECT 0.000000 537.000000 5.260000 538.080000 ;
      RECT 0.000000 536.580000 548.960000 537.000000 ;
      RECT 0.000000 535.360000 550.160000 536.580000 ;
      RECT 547.900000 535.120000 550.160000 535.360000 ;
      RECT 547.900000 534.280000 548.960000 535.120000 ;
      RECT 506.620000 534.280000 545.300000 535.360000 ;
      RECT 461.620000 534.280000 504.820000 535.360000 ;
      RECT 416.620000 534.280000 459.820000 535.360000 ;
      RECT 371.620000 534.280000 414.820000 535.360000 ;
      RECT 326.620000 534.280000 369.820000 535.360000 ;
      RECT 281.620000 534.280000 324.820000 535.360000 ;
      RECT 236.620000 534.280000 279.820000 535.360000 ;
      RECT 191.620000 534.280000 234.820000 535.360000 ;
      RECT 146.620000 534.280000 189.820000 535.360000 ;
      RECT 101.620000 534.280000 144.820000 535.360000 ;
      RECT 56.620000 534.280000 99.820000 535.360000 ;
      RECT 11.620000 534.280000 54.820000 535.360000 ;
      RECT 4.860000 534.280000 9.655000 535.360000 ;
      RECT 0.000000 534.280000 2.260000 535.360000 ;
      RECT 0.000000 534.140000 548.960000 534.280000 ;
      RECT 0.000000 532.680000 550.160000 534.140000 ;
      RECT 0.000000 532.640000 548.960000 532.680000 ;
      RECT 544.900000 531.700000 548.960000 532.640000 ;
      RECT 544.900000 531.560000 550.160000 531.700000 ;
      RECT 508.620000 531.560000 542.300000 532.640000 ;
      RECT 463.620000 531.560000 506.820000 532.640000 ;
      RECT 418.620000 531.560000 461.820000 532.640000 ;
      RECT 373.620000 531.560000 416.820000 532.640000 ;
      RECT 328.620000 531.560000 371.820000 532.640000 ;
      RECT 283.620000 531.560000 326.820000 532.640000 ;
      RECT 238.620000 531.560000 281.820000 532.640000 ;
      RECT 193.620000 531.560000 236.820000 532.640000 ;
      RECT 148.620000 531.560000 191.820000 532.640000 ;
      RECT 103.620000 531.560000 146.820000 532.640000 ;
      RECT 58.620000 531.560000 101.820000 532.640000 ;
      RECT 13.620000 531.560000 56.820000 532.640000 ;
      RECT 7.860000 531.560000 11.820000 532.640000 ;
      RECT 0.000000 531.560000 5.260000 532.640000 ;
      RECT 0.000000 530.240000 550.160000 531.560000 ;
      RECT 0.000000 529.920000 548.960000 530.240000 ;
      RECT 547.900000 529.260000 548.960000 529.920000 ;
      RECT 547.900000 528.840000 550.160000 529.260000 ;
      RECT 506.620000 528.840000 545.300000 529.920000 ;
      RECT 461.620000 528.840000 504.820000 529.920000 ;
      RECT 416.620000 528.840000 459.820000 529.920000 ;
      RECT 371.620000 528.840000 414.820000 529.920000 ;
      RECT 326.620000 528.840000 369.820000 529.920000 ;
      RECT 281.620000 528.840000 324.820000 529.920000 ;
      RECT 236.620000 528.840000 279.820000 529.920000 ;
      RECT 191.620000 528.840000 234.820000 529.920000 ;
      RECT 146.620000 528.840000 189.820000 529.920000 ;
      RECT 101.620000 528.840000 144.820000 529.920000 ;
      RECT 56.620000 528.840000 99.820000 529.920000 ;
      RECT 11.620000 528.840000 54.820000 529.920000 ;
      RECT 4.860000 528.840000 9.655000 529.920000 ;
      RECT 0.000000 528.840000 2.260000 529.920000 ;
      RECT 0.000000 528.410000 550.160000 528.840000 ;
      RECT 0.000000 527.430000 548.960000 528.410000 ;
      RECT 0.000000 527.200000 550.160000 527.430000 ;
      RECT 544.900000 526.120000 550.160000 527.200000 ;
      RECT 508.620000 526.120000 542.300000 527.200000 ;
      RECT 463.620000 526.120000 506.820000 527.200000 ;
      RECT 418.620000 526.120000 461.820000 527.200000 ;
      RECT 373.620000 526.120000 416.820000 527.200000 ;
      RECT 328.620000 526.120000 371.820000 527.200000 ;
      RECT 283.620000 526.120000 326.820000 527.200000 ;
      RECT 238.620000 526.120000 281.820000 527.200000 ;
      RECT 193.620000 526.120000 236.820000 527.200000 ;
      RECT 148.620000 526.120000 191.820000 527.200000 ;
      RECT 103.620000 526.120000 146.820000 527.200000 ;
      RECT 58.620000 526.120000 101.820000 527.200000 ;
      RECT 13.620000 526.120000 56.820000 527.200000 ;
      RECT 7.860000 526.120000 11.820000 527.200000 ;
      RECT 0.000000 526.120000 5.260000 527.200000 ;
      RECT 0.000000 525.970000 550.160000 526.120000 ;
      RECT 0.000000 524.990000 548.960000 525.970000 ;
      RECT 0.000000 524.480000 550.160000 524.990000 ;
      RECT 547.900000 523.530000 550.160000 524.480000 ;
      RECT 547.900000 523.400000 548.960000 523.530000 ;
      RECT 506.620000 523.400000 545.300000 524.480000 ;
      RECT 461.620000 523.400000 504.820000 524.480000 ;
      RECT 416.620000 523.400000 459.820000 524.480000 ;
      RECT 371.620000 523.400000 414.820000 524.480000 ;
      RECT 326.620000 523.400000 369.820000 524.480000 ;
      RECT 281.620000 523.400000 324.820000 524.480000 ;
      RECT 236.620000 523.400000 279.820000 524.480000 ;
      RECT 191.620000 523.400000 234.820000 524.480000 ;
      RECT 146.620000 523.400000 189.820000 524.480000 ;
      RECT 101.620000 523.400000 144.820000 524.480000 ;
      RECT 56.620000 523.400000 99.820000 524.480000 ;
      RECT 11.620000 523.400000 54.820000 524.480000 ;
      RECT 4.860000 523.400000 9.655000 524.480000 ;
      RECT 0.000000 523.400000 2.260000 524.480000 ;
      RECT 0.000000 522.550000 548.960000 523.400000 ;
      RECT 0.000000 521.760000 550.160000 522.550000 ;
      RECT 544.900000 521.090000 550.160000 521.760000 ;
      RECT 544.900000 520.680000 548.960000 521.090000 ;
      RECT 508.620000 520.680000 542.300000 521.760000 ;
      RECT 463.620000 520.680000 506.820000 521.760000 ;
      RECT 418.620000 520.680000 461.820000 521.760000 ;
      RECT 373.620000 520.680000 416.820000 521.760000 ;
      RECT 328.620000 520.680000 371.820000 521.760000 ;
      RECT 283.620000 520.680000 326.820000 521.760000 ;
      RECT 238.620000 520.680000 281.820000 521.760000 ;
      RECT 193.620000 520.680000 236.820000 521.760000 ;
      RECT 148.620000 520.680000 191.820000 521.760000 ;
      RECT 103.620000 520.680000 146.820000 521.760000 ;
      RECT 58.620000 520.680000 101.820000 521.760000 ;
      RECT 13.620000 520.680000 56.820000 521.760000 ;
      RECT 7.860000 520.680000 11.820000 521.760000 ;
      RECT 0.000000 520.680000 5.260000 521.760000 ;
      RECT 0.000000 520.110000 548.960000 520.680000 ;
      RECT 0.000000 519.260000 550.160000 520.110000 ;
      RECT 0.000000 519.040000 548.960000 519.260000 ;
      RECT 547.900000 518.280000 548.960000 519.040000 ;
      RECT 547.900000 517.960000 550.160000 518.280000 ;
      RECT 506.620000 517.960000 545.300000 519.040000 ;
      RECT 461.620000 517.960000 504.820000 519.040000 ;
      RECT 416.620000 517.960000 459.820000 519.040000 ;
      RECT 371.620000 517.960000 414.820000 519.040000 ;
      RECT 326.620000 517.960000 369.820000 519.040000 ;
      RECT 281.620000 517.960000 324.820000 519.040000 ;
      RECT 236.620000 517.960000 279.820000 519.040000 ;
      RECT 191.620000 517.960000 234.820000 519.040000 ;
      RECT 146.620000 517.960000 189.820000 519.040000 ;
      RECT 101.620000 517.960000 144.820000 519.040000 ;
      RECT 56.620000 517.960000 99.820000 519.040000 ;
      RECT 11.620000 517.960000 54.820000 519.040000 ;
      RECT 4.860000 517.960000 9.655000 519.040000 ;
      RECT 0.000000 517.960000 2.260000 519.040000 ;
      RECT 0.000000 516.820000 550.160000 517.960000 ;
      RECT 0.000000 516.320000 548.960000 516.820000 ;
      RECT 544.900000 515.840000 548.960000 516.320000 ;
      RECT 544.900000 515.240000 550.160000 515.840000 ;
      RECT 508.620000 515.240000 542.300000 516.320000 ;
      RECT 463.620000 515.240000 506.820000 516.320000 ;
      RECT 418.620000 515.240000 461.820000 516.320000 ;
      RECT 373.620000 515.240000 416.820000 516.320000 ;
      RECT 328.620000 515.240000 371.820000 516.320000 ;
      RECT 283.620000 515.240000 326.820000 516.320000 ;
      RECT 238.620000 515.240000 281.820000 516.320000 ;
      RECT 193.620000 515.240000 236.820000 516.320000 ;
      RECT 148.620000 515.240000 191.820000 516.320000 ;
      RECT 103.620000 515.240000 146.820000 516.320000 ;
      RECT 58.620000 515.240000 101.820000 516.320000 ;
      RECT 13.620000 515.240000 56.820000 516.320000 ;
      RECT 7.860000 515.240000 11.820000 516.320000 ;
      RECT 0.000000 515.240000 5.260000 516.320000 ;
      RECT 0.000000 514.380000 550.160000 515.240000 ;
      RECT 0.000000 513.600000 548.960000 514.380000 ;
      RECT 547.900000 513.400000 548.960000 513.600000 ;
      RECT 547.900000 512.520000 550.160000 513.400000 ;
      RECT 506.620000 512.520000 545.300000 513.600000 ;
      RECT 461.620000 512.520000 504.820000 513.600000 ;
      RECT 416.620000 512.520000 459.820000 513.600000 ;
      RECT 371.620000 512.520000 414.820000 513.600000 ;
      RECT 326.620000 512.520000 369.820000 513.600000 ;
      RECT 281.620000 512.520000 324.820000 513.600000 ;
      RECT 236.620000 512.520000 279.820000 513.600000 ;
      RECT 191.620000 512.520000 234.820000 513.600000 ;
      RECT 146.620000 512.520000 189.820000 513.600000 ;
      RECT 101.620000 512.520000 144.820000 513.600000 ;
      RECT 56.620000 512.520000 99.820000 513.600000 ;
      RECT 11.620000 512.520000 54.820000 513.600000 ;
      RECT 4.860000 512.520000 9.655000 513.600000 ;
      RECT 0.000000 512.520000 2.260000 513.600000 ;
      RECT 0.000000 511.940000 550.160000 512.520000 ;
      RECT 0.000000 510.960000 548.960000 511.940000 ;
      RECT 0.000000 510.880000 550.160000 510.960000 ;
      RECT 544.900000 510.110000 550.160000 510.880000 ;
      RECT 544.900000 509.800000 548.960000 510.110000 ;
      RECT 508.620000 509.800000 542.300000 510.880000 ;
      RECT 463.620000 509.800000 506.820000 510.880000 ;
      RECT 418.620000 509.800000 461.820000 510.880000 ;
      RECT 373.620000 509.800000 416.820000 510.880000 ;
      RECT 328.620000 509.800000 371.820000 510.880000 ;
      RECT 283.620000 509.800000 326.820000 510.880000 ;
      RECT 238.620000 509.800000 281.820000 510.880000 ;
      RECT 193.620000 509.800000 236.820000 510.880000 ;
      RECT 148.620000 509.800000 191.820000 510.880000 ;
      RECT 103.620000 509.800000 146.820000 510.880000 ;
      RECT 58.620000 509.800000 101.820000 510.880000 ;
      RECT 13.620000 509.800000 56.820000 510.880000 ;
      RECT 7.860000 509.800000 11.820000 510.880000 ;
      RECT 0.000000 509.800000 5.260000 510.880000 ;
      RECT 0.000000 509.130000 548.960000 509.800000 ;
      RECT 0.000000 508.160000 550.160000 509.130000 ;
      RECT 547.900000 507.670000 550.160000 508.160000 ;
      RECT 547.900000 507.080000 548.960000 507.670000 ;
      RECT 506.620000 507.080000 545.300000 508.160000 ;
      RECT 461.620000 507.080000 504.820000 508.160000 ;
      RECT 416.620000 507.080000 459.820000 508.160000 ;
      RECT 371.620000 507.080000 414.820000 508.160000 ;
      RECT 326.620000 507.080000 369.820000 508.160000 ;
      RECT 281.620000 507.080000 324.820000 508.160000 ;
      RECT 236.620000 507.080000 279.820000 508.160000 ;
      RECT 191.620000 507.080000 234.820000 508.160000 ;
      RECT 146.620000 507.080000 189.820000 508.160000 ;
      RECT 101.620000 507.080000 144.820000 508.160000 ;
      RECT 56.620000 507.080000 99.820000 508.160000 ;
      RECT 11.620000 507.080000 54.820000 508.160000 ;
      RECT 4.860000 507.080000 9.655000 508.160000 ;
      RECT 0.000000 507.080000 2.260000 508.160000 ;
      RECT 0.000000 506.690000 548.960000 507.080000 ;
      RECT 0.000000 505.440000 550.160000 506.690000 ;
      RECT 544.900000 505.230000 550.160000 505.440000 ;
      RECT 544.900000 504.360000 548.960000 505.230000 ;
      RECT 508.620000 504.360000 542.300000 505.440000 ;
      RECT 463.620000 504.360000 506.820000 505.440000 ;
      RECT 418.620000 504.360000 461.820000 505.440000 ;
      RECT 373.620000 504.360000 416.820000 505.440000 ;
      RECT 328.620000 504.360000 371.820000 505.440000 ;
      RECT 283.620000 504.360000 326.820000 505.440000 ;
      RECT 238.620000 504.360000 281.820000 505.440000 ;
      RECT 193.620000 504.360000 236.820000 505.440000 ;
      RECT 148.620000 504.360000 191.820000 505.440000 ;
      RECT 103.620000 504.360000 146.820000 505.440000 ;
      RECT 58.620000 504.360000 101.820000 505.440000 ;
      RECT 13.620000 504.360000 56.820000 505.440000 ;
      RECT 7.860000 504.360000 11.820000 505.440000 ;
      RECT 0.000000 504.360000 5.260000 505.440000 ;
      RECT 0.000000 504.250000 548.960000 504.360000 ;
      RECT 0.000000 502.790000 550.160000 504.250000 ;
      RECT 0.000000 502.720000 548.960000 502.790000 ;
      RECT 547.900000 501.810000 548.960000 502.720000 ;
      RECT 547.900000 501.640000 550.160000 501.810000 ;
      RECT 506.620000 501.640000 545.300000 502.720000 ;
      RECT 461.620000 501.640000 504.820000 502.720000 ;
      RECT 416.620000 501.640000 459.820000 502.720000 ;
      RECT 371.620000 501.640000 414.820000 502.720000 ;
      RECT 326.620000 501.640000 369.820000 502.720000 ;
      RECT 281.620000 501.640000 324.820000 502.720000 ;
      RECT 236.620000 501.640000 279.820000 502.720000 ;
      RECT 191.620000 501.640000 234.820000 502.720000 ;
      RECT 146.620000 501.640000 189.820000 502.720000 ;
      RECT 101.620000 501.640000 144.820000 502.720000 ;
      RECT 56.620000 501.640000 99.820000 502.720000 ;
      RECT 11.620000 501.640000 54.820000 502.720000 ;
      RECT 4.860000 501.640000 9.655000 502.720000 ;
      RECT 0.000000 501.640000 2.260000 502.720000 ;
      RECT 0.000000 500.960000 550.160000 501.640000 ;
      RECT 0.000000 500.000000 548.960000 500.960000 ;
      RECT 544.900000 499.980000 548.960000 500.000000 ;
      RECT 544.900000 498.920000 550.160000 499.980000 ;
      RECT 508.620000 498.920000 542.300000 500.000000 ;
      RECT 463.620000 498.920000 506.820000 500.000000 ;
      RECT 418.620000 498.920000 461.820000 500.000000 ;
      RECT 373.620000 498.920000 416.820000 500.000000 ;
      RECT 328.620000 498.920000 371.820000 500.000000 ;
      RECT 283.620000 498.920000 326.820000 500.000000 ;
      RECT 238.620000 498.920000 281.820000 500.000000 ;
      RECT 193.620000 498.920000 236.820000 500.000000 ;
      RECT 148.620000 498.920000 191.820000 500.000000 ;
      RECT 103.620000 498.920000 146.820000 500.000000 ;
      RECT 58.620000 498.920000 101.820000 500.000000 ;
      RECT 13.620000 498.920000 56.820000 500.000000 ;
      RECT 7.860000 498.920000 11.820000 500.000000 ;
      RECT 0.000000 498.920000 5.260000 500.000000 ;
      RECT 0.000000 498.520000 550.160000 498.920000 ;
      RECT 0.000000 497.540000 548.960000 498.520000 ;
      RECT 0.000000 497.280000 550.160000 497.540000 ;
      RECT 547.900000 496.200000 550.160000 497.280000 ;
      RECT 506.620000 496.200000 545.300000 497.280000 ;
      RECT 461.620000 496.200000 504.820000 497.280000 ;
      RECT 416.620000 496.200000 459.820000 497.280000 ;
      RECT 371.620000 496.200000 414.820000 497.280000 ;
      RECT 326.620000 496.200000 369.820000 497.280000 ;
      RECT 281.620000 496.200000 324.820000 497.280000 ;
      RECT 236.620000 496.200000 279.820000 497.280000 ;
      RECT 191.620000 496.200000 234.820000 497.280000 ;
      RECT 146.620000 496.200000 189.820000 497.280000 ;
      RECT 101.620000 496.200000 144.820000 497.280000 ;
      RECT 56.620000 496.200000 99.820000 497.280000 ;
      RECT 11.620000 496.200000 54.820000 497.280000 ;
      RECT 4.860000 496.200000 9.655000 497.280000 ;
      RECT 0.000000 496.200000 2.260000 497.280000 ;
      RECT 0.000000 496.080000 550.160000 496.200000 ;
      RECT 0.000000 495.100000 548.960000 496.080000 ;
      RECT 0.000000 494.560000 550.160000 495.100000 ;
      RECT 544.900000 493.640000 550.160000 494.560000 ;
      RECT 544.900000 493.480000 548.960000 493.640000 ;
      RECT 508.620000 493.480000 542.300000 494.560000 ;
      RECT 463.620000 493.480000 506.820000 494.560000 ;
      RECT 418.620000 493.480000 461.820000 494.560000 ;
      RECT 373.620000 493.480000 416.820000 494.560000 ;
      RECT 328.620000 493.480000 371.820000 494.560000 ;
      RECT 283.620000 493.480000 326.820000 494.560000 ;
      RECT 238.620000 493.480000 281.820000 494.560000 ;
      RECT 193.620000 493.480000 236.820000 494.560000 ;
      RECT 148.620000 493.480000 191.820000 494.560000 ;
      RECT 103.620000 493.480000 146.820000 494.560000 ;
      RECT 58.620000 493.480000 101.820000 494.560000 ;
      RECT 13.620000 493.480000 56.820000 494.560000 ;
      RECT 7.860000 493.480000 11.820000 494.560000 ;
      RECT 0.000000 493.480000 5.260000 494.560000 ;
      RECT 0.000000 492.660000 548.960000 493.480000 ;
      RECT 0.000000 491.840000 550.160000 492.660000 ;
      RECT 547.900000 491.810000 550.160000 491.840000 ;
      RECT 547.900000 490.830000 548.960000 491.810000 ;
      RECT 547.900000 490.760000 550.160000 490.830000 ;
      RECT 506.620000 490.760000 545.300000 491.840000 ;
      RECT 461.620000 490.760000 504.820000 491.840000 ;
      RECT 416.620000 490.760000 459.820000 491.840000 ;
      RECT 371.620000 490.760000 414.820000 491.840000 ;
      RECT 326.620000 490.760000 369.820000 491.840000 ;
      RECT 281.620000 490.760000 324.820000 491.840000 ;
      RECT 236.620000 490.760000 279.820000 491.840000 ;
      RECT 191.620000 490.760000 234.820000 491.840000 ;
      RECT 146.620000 490.760000 189.820000 491.840000 ;
      RECT 101.620000 490.760000 144.820000 491.840000 ;
      RECT 56.620000 490.760000 99.820000 491.840000 ;
      RECT 11.620000 490.760000 54.820000 491.840000 ;
      RECT 4.860000 490.760000 9.655000 491.840000 ;
      RECT 0.000000 490.760000 2.260000 491.840000 ;
      RECT 0.000000 489.370000 550.160000 490.760000 ;
      RECT 0.000000 489.120000 548.960000 489.370000 ;
      RECT 544.900000 488.390000 548.960000 489.120000 ;
      RECT 544.900000 488.040000 550.160000 488.390000 ;
      RECT 508.620000 488.040000 542.300000 489.120000 ;
      RECT 463.620000 488.040000 506.820000 489.120000 ;
      RECT 418.620000 488.040000 461.820000 489.120000 ;
      RECT 373.620000 488.040000 416.820000 489.120000 ;
      RECT 328.620000 488.040000 371.820000 489.120000 ;
      RECT 283.620000 488.040000 326.820000 489.120000 ;
      RECT 238.620000 488.040000 281.820000 489.120000 ;
      RECT 193.620000 488.040000 236.820000 489.120000 ;
      RECT 148.620000 488.040000 191.820000 489.120000 ;
      RECT 103.620000 488.040000 146.820000 489.120000 ;
      RECT 58.620000 488.040000 101.820000 489.120000 ;
      RECT 13.620000 488.040000 56.820000 489.120000 ;
      RECT 7.860000 488.040000 11.820000 489.120000 ;
      RECT 0.000000 488.040000 5.260000 489.120000 ;
      RECT 0.000000 486.930000 550.160000 488.040000 ;
      RECT 0.000000 486.400000 548.960000 486.930000 ;
      RECT 547.900000 485.950000 548.960000 486.400000 ;
      RECT 547.900000 485.320000 550.160000 485.950000 ;
      RECT 506.620000 485.320000 545.300000 486.400000 ;
      RECT 461.620000 485.320000 504.820000 486.400000 ;
      RECT 416.620000 485.320000 459.820000 486.400000 ;
      RECT 371.620000 485.320000 414.820000 486.400000 ;
      RECT 326.620000 485.320000 369.820000 486.400000 ;
      RECT 281.620000 485.320000 324.820000 486.400000 ;
      RECT 236.620000 485.320000 279.820000 486.400000 ;
      RECT 191.620000 485.320000 234.820000 486.400000 ;
      RECT 146.620000 485.320000 189.820000 486.400000 ;
      RECT 101.620000 485.320000 144.820000 486.400000 ;
      RECT 56.620000 485.320000 99.820000 486.400000 ;
      RECT 11.620000 485.320000 54.820000 486.400000 ;
      RECT 4.860000 485.320000 9.655000 486.400000 ;
      RECT 0.000000 485.320000 2.260000 486.400000 ;
      RECT 0.000000 484.490000 550.160000 485.320000 ;
      RECT 0.000000 483.680000 548.960000 484.490000 ;
      RECT 544.900000 483.510000 548.960000 483.680000 ;
      RECT 544.900000 482.660000 550.160000 483.510000 ;
      RECT 544.900000 482.600000 548.960000 482.660000 ;
      RECT 508.620000 482.600000 542.300000 483.680000 ;
      RECT 463.620000 482.600000 506.820000 483.680000 ;
      RECT 418.620000 482.600000 461.820000 483.680000 ;
      RECT 373.620000 482.600000 416.820000 483.680000 ;
      RECT 328.620000 482.600000 371.820000 483.680000 ;
      RECT 283.620000 482.600000 326.820000 483.680000 ;
      RECT 238.620000 482.600000 281.820000 483.680000 ;
      RECT 193.620000 482.600000 236.820000 483.680000 ;
      RECT 148.620000 482.600000 191.820000 483.680000 ;
      RECT 103.620000 482.600000 146.820000 483.680000 ;
      RECT 58.620000 482.600000 101.820000 483.680000 ;
      RECT 13.620000 482.600000 56.820000 483.680000 ;
      RECT 7.860000 482.600000 11.820000 483.680000 ;
      RECT 0.000000 482.600000 5.260000 483.680000 ;
      RECT 0.000000 481.680000 548.960000 482.600000 ;
      RECT 0.000000 480.960000 550.160000 481.680000 ;
      RECT 547.900000 480.220000 550.160000 480.960000 ;
      RECT 547.900000 479.880000 548.960000 480.220000 ;
      RECT 506.620000 479.880000 545.300000 480.960000 ;
      RECT 461.620000 479.880000 504.820000 480.960000 ;
      RECT 416.620000 479.880000 459.820000 480.960000 ;
      RECT 371.620000 479.880000 414.820000 480.960000 ;
      RECT 326.620000 479.880000 369.820000 480.960000 ;
      RECT 281.620000 479.880000 324.820000 480.960000 ;
      RECT 236.620000 479.880000 279.820000 480.960000 ;
      RECT 191.620000 479.880000 234.820000 480.960000 ;
      RECT 146.620000 479.880000 189.820000 480.960000 ;
      RECT 101.620000 479.880000 144.820000 480.960000 ;
      RECT 56.620000 479.880000 99.820000 480.960000 ;
      RECT 11.620000 479.880000 54.820000 480.960000 ;
      RECT 4.860000 479.880000 9.655000 480.960000 ;
      RECT 0.000000 479.880000 2.260000 480.960000 ;
      RECT 0.000000 479.240000 548.960000 479.880000 ;
      RECT 0.000000 478.240000 550.160000 479.240000 ;
      RECT 544.900000 477.780000 550.160000 478.240000 ;
      RECT 544.900000 477.160000 548.960000 477.780000 ;
      RECT 508.620000 477.160000 542.300000 478.240000 ;
      RECT 463.620000 477.160000 506.820000 478.240000 ;
      RECT 418.620000 477.160000 461.820000 478.240000 ;
      RECT 373.620000 477.160000 416.820000 478.240000 ;
      RECT 328.620000 477.160000 371.820000 478.240000 ;
      RECT 283.620000 477.160000 326.820000 478.240000 ;
      RECT 238.620000 477.160000 281.820000 478.240000 ;
      RECT 193.620000 477.160000 236.820000 478.240000 ;
      RECT 148.620000 477.160000 191.820000 478.240000 ;
      RECT 103.620000 477.160000 146.820000 478.240000 ;
      RECT 58.620000 477.160000 101.820000 478.240000 ;
      RECT 13.620000 477.160000 56.820000 478.240000 ;
      RECT 7.860000 477.160000 11.820000 478.240000 ;
      RECT 0.000000 477.160000 5.260000 478.240000 ;
      RECT 0.000000 476.800000 548.960000 477.160000 ;
      RECT 0.000000 475.520000 550.160000 476.800000 ;
      RECT 547.900000 475.340000 550.160000 475.520000 ;
      RECT 547.900000 474.440000 548.960000 475.340000 ;
      RECT 506.620000 474.440000 545.300000 475.520000 ;
      RECT 461.620000 474.440000 504.820000 475.520000 ;
      RECT 416.620000 474.440000 459.820000 475.520000 ;
      RECT 371.620000 474.440000 414.820000 475.520000 ;
      RECT 326.620000 474.440000 369.820000 475.520000 ;
      RECT 281.620000 474.440000 324.820000 475.520000 ;
      RECT 236.620000 474.440000 279.820000 475.520000 ;
      RECT 191.620000 474.440000 234.820000 475.520000 ;
      RECT 146.620000 474.440000 189.820000 475.520000 ;
      RECT 101.620000 474.440000 144.820000 475.520000 ;
      RECT 56.620000 474.440000 99.820000 475.520000 ;
      RECT 11.620000 474.440000 54.820000 475.520000 ;
      RECT 4.860000 474.440000 9.655000 475.520000 ;
      RECT 0.000000 474.440000 2.260000 475.520000 ;
      RECT 0.000000 474.360000 548.960000 474.440000 ;
      RECT 0.000000 473.510000 550.160000 474.360000 ;
      RECT 0.000000 472.800000 548.960000 473.510000 ;
      RECT 544.900000 472.530000 548.960000 472.800000 ;
      RECT 544.900000 471.720000 550.160000 472.530000 ;
      RECT 508.620000 471.720000 542.300000 472.800000 ;
      RECT 463.620000 471.720000 506.820000 472.800000 ;
      RECT 418.620000 471.720000 461.820000 472.800000 ;
      RECT 373.620000 471.720000 416.820000 472.800000 ;
      RECT 328.620000 471.720000 371.820000 472.800000 ;
      RECT 283.620000 471.720000 326.820000 472.800000 ;
      RECT 238.620000 471.720000 281.820000 472.800000 ;
      RECT 193.620000 471.720000 236.820000 472.800000 ;
      RECT 148.620000 471.720000 191.820000 472.800000 ;
      RECT 103.620000 471.720000 146.820000 472.800000 ;
      RECT 58.620000 471.720000 101.820000 472.800000 ;
      RECT 13.620000 471.720000 56.820000 472.800000 ;
      RECT 7.860000 471.720000 11.820000 472.800000 ;
      RECT 0.000000 471.720000 5.260000 472.800000 ;
      RECT 0.000000 471.070000 550.160000 471.720000 ;
      RECT 0.000000 470.090000 548.960000 471.070000 ;
      RECT 0.000000 470.080000 550.160000 470.090000 ;
      RECT 547.900000 469.000000 550.160000 470.080000 ;
      RECT 506.620000 469.000000 545.300000 470.080000 ;
      RECT 461.620000 469.000000 504.820000 470.080000 ;
      RECT 416.620000 469.000000 459.820000 470.080000 ;
      RECT 371.620000 469.000000 414.820000 470.080000 ;
      RECT 326.620000 469.000000 369.820000 470.080000 ;
      RECT 281.620000 469.000000 324.820000 470.080000 ;
      RECT 236.620000 469.000000 279.820000 470.080000 ;
      RECT 191.620000 469.000000 234.820000 470.080000 ;
      RECT 146.620000 469.000000 189.820000 470.080000 ;
      RECT 101.620000 469.000000 144.820000 470.080000 ;
      RECT 56.620000 469.000000 99.820000 470.080000 ;
      RECT 11.620000 469.000000 54.820000 470.080000 ;
      RECT 4.860000 469.000000 9.655000 470.080000 ;
      RECT 0.000000 469.000000 2.260000 470.080000 ;
      RECT 0.000000 468.630000 550.160000 469.000000 ;
      RECT 0.000000 467.650000 548.960000 468.630000 ;
      RECT 0.000000 467.360000 550.160000 467.650000 ;
      RECT 544.900000 466.280000 550.160000 467.360000 ;
      RECT 508.620000 466.280000 542.300000 467.360000 ;
      RECT 463.620000 466.280000 506.820000 467.360000 ;
      RECT 418.620000 466.280000 461.820000 467.360000 ;
      RECT 373.620000 466.280000 416.820000 467.360000 ;
      RECT 328.620000 466.280000 371.820000 467.360000 ;
      RECT 283.620000 466.280000 326.820000 467.360000 ;
      RECT 238.620000 466.280000 281.820000 467.360000 ;
      RECT 193.620000 466.280000 236.820000 467.360000 ;
      RECT 148.620000 466.280000 191.820000 467.360000 ;
      RECT 103.620000 466.280000 146.820000 467.360000 ;
      RECT 58.620000 466.280000 101.820000 467.360000 ;
      RECT 13.620000 466.280000 56.820000 467.360000 ;
      RECT 7.860000 466.280000 11.820000 467.360000 ;
      RECT 0.000000 466.280000 5.260000 467.360000 ;
      RECT 0.000000 466.190000 550.160000 466.280000 ;
      RECT 0.000000 465.210000 548.960000 466.190000 ;
      RECT 0.000000 464.640000 550.160000 465.210000 ;
      RECT 547.900000 463.750000 550.160000 464.640000 ;
      RECT 547.900000 463.560000 548.960000 463.750000 ;
      RECT 506.620000 463.560000 545.300000 464.640000 ;
      RECT 461.620000 463.560000 504.820000 464.640000 ;
      RECT 416.620000 463.560000 459.820000 464.640000 ;
      RECT 371.620000 463.560000 414.820000 464.640000 ;
      RECT 326.620000 463.560000 369.820000 464.640000 ;
      RECT 281.620000 463.560000 324.820000 464.640000 ;
      RECT 236.620000 463.560000 279.820000 464.640000 ;
      RECT 191.620000 463.560000 234.820000 464.640000 ;
      RECT 146.620000 463.560000 189.820000 464.640000 ;
      RECT 101.620000 463.560000 144.820000 464.640000 ;
      RECT 56.620000 463.560000 99.820000 464.640000 ;
      RECT 11.620000 463.560000 54.820000 464.640000 ;
      RECT 4.860000 463.560000 9.655000 464.640000 ;
      RECT 0.000000 463.560000 2.260000 464.640000 ;
      RECT 0.000000 462.770000 548.960000 463.560000 ;
      RECT 0.000000 461.920000 550.160000 462.770000 ;
      RECT 544.900000 460.940000 548.960000 461.920000 ;
      RECT 544.900000 460.840000 550.160000 460.940000 ;
      RECT 508.620000 460.840000 542.300000 461.920000 ;
      RECT 463.620000 460.840000 506.820000 461.920000 ;
      RECT 418.620000 460.840000 461.820000 461.920000 ;
      RECT 373.620000 460.840000 416.820000 461.920000 ;
      RECT 328.620000 460.840000 371.820000 461.920000 ;
      RECT 283.620000 460.840000 326.820000 461.920000 ;
      RECT 238.620000 460.840000 281.820000 461.920000 ;
      RECT 193.620000 460.840000 236.820000 461.920000 ;
      RECT 148.620000 460.840000 191.820000 461.920000 ;
      RECT 103.620000 460.840000 146.820000 461.920000 ;
      RECT 58.620000 460.840000 101.820000 461.920000 ;
      RECT 13.620000 460.840000 56.820000 461.920000 ;
      RECT 7.860000 460.840000 11.820000 461.920000 ;
      RECT 0.000000 460.840000 5.260000 461.920000 ;
      RECT 0.000000 459.480000 550.160000 460.840000 ;
      RECT 0.000000 459.200000 548.960000 459.480000 ;
      RECT 547.900000 458.500000 548.960000 459.200000 ;
      RECT 547.900000 458.120000 550.160000 458.500000 ;
      RECT 506.620000 458.120000 545.300000 459.200000 ;
      RECT 461.620000 458.120000 504.820000 459.200000 ;
      RECT 416.620000 458.120000 459.820000 459.200000 ;
      RECT 371.620000 458.120000 414.820000 459.200000 ;
      RECT 326.620000 458.120000 369.820000 459.200000 ;
      RECT 281.620000 458.120000 324.820000 459.200000 ;
      RECT 236.620000 458.120000 279.820000 459.200000 ;
      RECT 191.620000 458.120000 234.820000 459.200000 ;
      RECT 146.620000 458.120000 189.820000 459.200000 ;
      RECT 101.620000 458.120000 144.820000 459.200000 ;
      RECT 56.620000 458.120000 99.820000 459.200000 ;
      RECT 11.620000 458.120000 54.820000 459.200000 ;
      RECT 4.860000 458.120000 9.655000 459.200000 ;
      RECT 0.000000 458.120000 2.260000 459.200000 ;
      RECT 0.000000 457.040000 550.160000 458.120000 ;
      RECT 0.000000 456.480000 548.960000 457.040000 ;
      RECT 544.900000 456.060000 548.960000 456.480000 ;
      RECT 544.900000 455.400000 550.160000 456.060000 ;
      RECT 508.620000 455.400000 542.300000 456.480000 ;
      RECT 463.620000 455.400000 506.820000 456.480000 ;
      RECT 418.620000 455.400000 461.820000 456.480000 ;
      RECT 373.620000 455.400000 416.820000 456.480000 ;
      RECT 328.620000 455.400000 371.820000 456.480000 ;
      RECT 283.620000 455.400000 326.820000 456.480000 ;
      RECT 238.620000 455.400000 281.820000 456.480000 ;
      RECT 193.620000 455.400000 236.820000 456.480000 ;
      RECT 148.620000 455.400000 191.820000 456.480000 ;
      RECT 103.620000 455.400000 146.820000 456.480000 ;
      RECT 58.620000 455.400000 101.820000 456.480000 ;
      RECT 13.620000 455.400000 56.820000 456.480000 ;
      RECT 7.860000 455.400000 11.820000 456.480000 ;
      RECT 0.000000 455.400000 5.260000 456.480000 ;
      RECT 0.000000 454.600000 550.160000 455.400000 ;
      RECT 0.000000 453.760000 548.960000 454.600000 ;
      RECT 547.900000 453.620000 548.960000 453.760000 ;
      RECT 547.900000 452.770000 550.160000 453.620000 ;
      RECT 547.900000 452.680000 548.960000 452.770000 ;
      RECT 506.620000 452.680000 545.300000 453.760000 ;
      RECT 461.620000 452.680000 504.820000 453.760000 ;
      RECT 416.620000 452.680000 459.820000 453.760000 ;
      RECT 371.620000 452.680000 414.820000 453.760000 ;
      RECT 326.620000 452.680000 369.820000 453.760000 ;
      RECT 281.620000 452.680000 324.820000 453.760000 ;
      RECT 236.620000 452.680000 279.820000 453.760000 ;
      RECT 191.620000 452.680000 234.820000 453.760000 ;
      RECT 146.620000 452.680000 189.820000 453.760000 ;
      RECT 101.620000 452.680000 144.820000 453.760000 ;
      RECT 56.620000 452.680000 99.820000 453.760000 ;
      RECT 11.620000 452.680000 54.820000 453.760000 ;
      RECT 4.860000 452.680000 9.655000 453.760000 ;
      RECT 0.000000 452.680000 2.260000 453.760000 ;
      RECT 0.000000 451.790000 548.960000 452.680000 ;
      RECT 0.000000 451.040000 550.160000 451.790000 ;
      RECT 544.900000 450.330000 550.160000 451.040000 ;
      RECT 544.900000 449.960000 548.960000 450.330000 ;
      RECT 508.620000 449.960000 542.300000 451.040000 ;
      RECT 463.620000 449.960000 506.820000 451.040000 ;
      RECT 418.620000 449.960000 461.820000 451.040000 ;
      RECT 373.620000 449.960000 416.820000 451.040000 ;
      RECT 328.620000 449.960000 371.820000 451.040000 ;
      RECT 283.620000 449.960000 326.820000 451.040000 ;
      RECT 238.620000 449.960000 281.820000 451.040000 ;
      RECT 193.620000 449.960000 236.820000 451.040000 ;
      RECT 148.620000 449.960000 191.820000 451.040000 ;
      RECT 103.620000 449.960000 146.820000 451.040000 ;
      RECT 58.620000 449.960000 101.820000 451.040000 ;
      RECT 13.620000 449.960000 56.820000 451.040000 ;
      RECT 7.860000 449.960000 11.820000 451.040000 ;
      RECT 0.000000 449.960000 5.260000 451.040000 ;
      RECT 0.000000 449.350000 548.960000 449.960000 ;
      RECT 0.000000 448.320000 550.160000 449.350000 ;
      RECT 547.900000 447.890000 550.160000 448.320000 ;
      RECT 547.900000 447.240000 548.960000 447.890000 ;
      RECT 506.620000 447.240000 545.300000 448.320000 ;
      RECT 461.620000 447.240000 504.820000 448.320000 ;
      RECT 416.620000 447.240000 459.820000 448.320000 ;
      RECT 371.620000 447.240000 414.820000 448.320000 ;
      RECT 326.620000 447.240000 369.820000 448.320000 ;
      RECT 281.620000 447.240000 324.820000 448.320000 ;
      RECT 236.620000 447.240000 279.820000 448.320000 ;
      RECT 191.620000 447.240000 234.820000 448.320000 ;
      RECT 146.620000 447.240000 189.820000 448.320000 ;
      RECT 101.620000 447.240000 144.820000 448.320000 ;
      RECT 56.620000 447.240000 99.820000 448.320000 ;
      RECT 11.620000 447.240000 54.820000 448.320000 ;
      RECT 4.860000 447.240000 9.655000 448.320000 ;
      RECT 0.000000 447.240000 2.260000 448.320000 ;
      RECT 0.000000 446.910000 548.960000 447.240000 ;
      RECT 0.000000 445.600000 550.160000 446.910000 ;
      RECT 544.900000 445.450000 550.160000 445.600000 ;
      RECT 544.900000 444.520000 548.960000 445.450000 ;
      RECT 508.620000 444.520000 542.300000 445.600000 ;
      RECT 463.620000 444.520000 506.820000 445.600000 ;
      RECT 418.620000 444.520000 461.820000 445.600000 ;
      RECT 373.620000 444.520000 416.820000 445.600000 ;
      RECT 328.620000 444.520000 371.820000 445.600000 ;
      RECT 283.620000 444.520000 326.820000 445.600000 ;
      RECT 238.620000 444.520000 281.820000 445.600000 ;
      RECT 193.620000 444.520000 236.820000 445.600000 ;
      RECT 148.620000 444.520000 191.820000 445.600000 ;
      RECT 103.620000 444.520000 146.820000 445.600000 ;
      RECT 58.620000 444.520000 101.820000 445.600000 ;
      RECT 13.620000 444.520000 56.820000 445.600000 ;
      RECT 7.860000 444.520000 11.820000 445.600000 ;
      RECT 0.000000 444.520000 5.260000 445.600000 ;
      RECT 0.000000 444.470000 548.960000 444.520000 ;
      RECT 0.000000 443.620000 550.160000 444.470000 ;
      RECT 0.000000 442.880000 548.960000 443.620000 ;
      RECT 547.900000 442.640000 548.960000 442.880000 ;
      RECT 547.900000 441.800000 550.160000 442.640000 ;
      RECT 506.620000 441.800000 545.300000 442.880000 ;
      RECT 461.620000 441.800000 504.820000 442.880000 ;
      RECT 416.620000 441.800000 459.820000 442.880000 ;
      RECT 371.620000 441.800000 414.820000 442.880000 ;
      RECT 326.620000 441.800000 369.820000 442.880000 ;
      RECT 281.620000 441.800000 324.820000 442.880000 ;
      RECT 236.620000 441.800000 279.820000 442.880000 ;
      RECT 191.620000 441.800000 234.820000 442.880000 ;
      RECT 146.620000 441.800000 189.820000 442.880000 ;
      RECT 101.620000 441.800000 144.820000 442.880000 ;
      RECT 56.620000 441.800000 99.820000 442.880000 ;
      RECT 11.620000 441.800000 54.820000 442.880000 ;
      RECT 4.860000 441.800000 9.655000 442.880000 ;
      RECT 0.000000 441.800000 2.260000 442.880000 ;
      RECT 0.000000 441.180000 550.160000 441.800000 ;
      RECT 0.000000 440.200000 548.960000 441.180000 ;
      RECT 0.000000 440.160000 550.160000 440.200000 ;
      RECT 544.900000 439.080000 550.160000 440.160000 ;
      RECT 508.620000 439.080000 542.300000 440.160000 ;
      RECT 463.620000 439.080000 506.820000 440.160000 ;
      RECT 418.620000 439.080000 461.820000 440.160000 ;
      RECT 373.620000 439.080000 416.820000 440.160000 ;
      RECT 328.620000 439.080000 371.820000 440.160000 ;
      RECT 283.620000 439.080000 326.820000 440.160000 ;
      RECT 238.620000 439.080000 281.820000 440.160000 ;
      RECT 193.620000 439.080000 236.820000 440.160000 ;
      RECT 148.620000 439.080000 191.820000 440.160000 ;
      RECT 103.620000 439.080000 146.820000 440.160000 ;
      RECT 58.620000 439.080000 101.820000 440.160000 ;
      RECT 13.620000 439.080000 56.820000 440.160000 ;
      RECT 7.860000 439.080000 11.820000 440.160000 ;
      RECT 0.000000 439.080000 5.260000 440.160000 ;
      RECT 0.000000 438.740000 550.160000 439.080000 ;
      RECT 0.000000 437.760000 548.960000 438.740000 ;
      RECT 0.000000 437.440000 550.160000 437.760000 ;
      RECT 547.900000 436.360000 550.160000 437.440000 ;
      RECT 506.620000 436.360000 545.300000 437.440000 ;
      RECT 461.620000 436.360000 504.820000 437.440000 ;
      RECT 416.620000 436.360000 459.820000 437.440000 ;
      RECT 371.620000 436.360000 414.820000 437.440000 ;
      RECT 326.620000 436.360000 369.820000 437.440000 ;
      RECT 281.620000 436.360000 324.820000 437.440000 ;
      RECT 236.620000 436.360000 279.820000 437.440000 ;
      RECT 191.620000 436.360000 234.820000 437.440000 ;
      RECT 146.620000 436.360000 189.820000 437.440000 ;
      RECT 101.620000 436.360000 144.820000 437.440000 ;
      RECT 56.620000 436.360000 99.820000 437.440000 ;
      RECT 11.620000 436.360000 54.820000 437.440000 ;
      RECT 4.860000 436.360000 9.655000 437.440000 ;
      RECT 0.000000 436.360000 2.260000 437.440000 ;
      RECT 0.000000 436.300000 550.160000 436.360000 ;
      RECT 0.000000 435.320000 548.960000 436.300000 ;
      RECT 0.000000 434.720000 550.160000 435.320000 ;
      RECT 544.900000 434.470000 550.160000 434.720000 ;
      RECT 544.900000 433.640000 548.960000 434.470000 ;
      RECT 508.620000 433.640000 542.300000 434.720000 ;
      RECT 463.620000 433.640000 506.820000 434.720000 ;
      RECT 418.620000 433.640000 461.820000 434.720000 ;
      RECT 373.620000 433.640000 416.820000 434.720000 ;
      RECT 328.620000 433.640000 371.820000 434.720000 ;
      RECT 283.620000 433.640000 326.820000 434.720000 ;
      RECT 238.620000 433.640000 281.820000 434.720000 ;
      RECT 193.620000 433.640000 236.820000 434.720000 ;
      RECT 148.620000 433.640000 191.820000 434.720000 ;
      RECT 103.620000 433.640000 146.820000 434.720000 ;
      RECT 58.620000 433.640000 101.820000 434.720000 ;
      RECT 13.620000 433.640000 56.820000 434.720000 ;
      RECT 7.860000 433.640000 11.820000 434.720000 ;
      RECT 0.000000 433.640000 5.260000 434.720000 ;
      RECT 0.000000 433.490000 548.960000 433.640000 ;
      RECT 0.000000 432.030000 550.160000 433.490000 ;
      RECT 0.000000 432.000000 548.960000 432.030000 ;
      RECT 547.900000 431.050000 548.960000 432.000000 ;
      RECT 547.900000 430.920000 550.160000 431.050000 ;
      RECT 506.620000 430.920000 545.300000 432.000000 ;
      RECT 461.620000 430.920000 504.820000 432.000000 ;
      RECT 416.620000 430.920000 459.820000 432.000000 ;
      RECT 371.620000 430.920000 414.820000 432.000000 ;
      RECT 326.620000 430.920000 369.820000 432.000000 ;
      RECT 281.620000 430.920000 324.820000 432.000000 ;
      RECT 236.620000 430.920000 279.820000 432.000000 ;
      RECT 191.620000 430.920000 234.820000 432.000000 ;
      RECT 146.620000 430.920000 189.820000 432.000000 ;
      RECT 101.620000 430.920000 144.820000 432.000000 ;
      RECT 56.620000 430.920000 99.820000 432.000000 ;
      RECT 11.620000 430.920000 54.820000 432.000000 ;
      RECT 4.860000 430.920000 9.655000 432.000000 ;
      RECT 0.000000 430.920000 2.260000 432.000000 ;
      RECT 0.000000 429.590000 550.160000 430.920000 ;
      RECT 0.000000 429.280000 548.960000 429.590000 ;
      RECT 544.900000 428.610000 548.960000 429.280000 ;
      RECT 544.900000 428.200000 550.160000 428.610000 ;
      RECT 508.620000 428.200000 542.300000 429.280000 ;
      RECT 463.620000 428.200000 506.820000 429.280000 ;
      RECT 418.620000 428.200000 461.820000 429.280000 ;
      RECT 373.620000 428.200000 416.820000 429.280000 ;
      RECT 328.620000 428.200000 371.820000 429.280000 ;
      RECT 283.620000 428.200000 326.820000 429.280000 ;
      RECT 238.620000 428.200000 281.820000 429.280000 ;
      RECT 193.620000 428.200000 236.820000 429.280000 ;
      RECT 148.620000 428.200000 191.820000 429.280000 ;
      RECT 103.620000 428.200000 146.820000 429.280000 ;
      RECT 58.620000 428.200000 101.820000 429.280000 ;
      RECT 13.620000 428.200000 56.820000 429.280000 ;
      RECT 7.860000 428.200000 11.820000 429.280000 ;
      RECT 0.000000 428.200000 5.260000 429.280000 ;
      RECT 0.000000 427.150000 550.160000 428.200000 ;
      RECT 0.000000 426.560000 548.960000 427.150000 ;
      RECT 547.900000 426.170000 548.960000 426.560000 ;
      RECT 547.900000 425.480000 550.160000 426.170000 ;
      RECT 506.620000 425.480000 545.300000 426.560000 ;
      RECT 461.620000 425.480000 504.820000 426.560000 ;
      RECT 416.620000 425.480000 459.820000 426.560000 ;
      RECT 371.620000 425.480000 414.820000 426.560000 ;
      RECT 326.620000 425.480000 369.820000 426.560000 ;
      RECT 281.620000 425.480000 324.820000 426.560000 ;
      RECT 236.620000 425.480000 279.820000 426.560000 ;
      RECT 191.620000 425.480000 234.820000 426.560000 ;
      RECT 146.620000 425.480000 189.820000 426.560000 ;
      RECT 101.620000 425.480000 144.820000 426.560000 ;
      RECT 56.620000 425.480000 99.820000 426.560000 ;
      RECT 11.620000 425.480000 54.820000 426.560000 ;
      RECT 4.860000 425.480000 9.655000 426.560000 ;
      RECT 0.000000 425.480000 2.260000 426.560000 ;
      RECT 0.000000 425.320000 550.160000 425.480000 ;
      RECT 0.000000 424.340000 548.960000 425.320000 ;
      RECT 0.000000 423.840000 550.160000 424.340000 ;
      RECT 544.900000 422.880000 550.160000 423.840000 ;
      RECT 544.900000 422.760000 548.960000 422.880000 ;
      RECT 508.620000 422.760000 542.300000 423.840000 ;
      RECT 463.620000 422.760000 506.820000 423.840000 ;
      RECT 418.620000 422.760000 461.820000 423.840000 ;
      RECT 373.620000 422.760000 416.820000 423.840000 ;
      RECT 328.620000 422.760000 371.820000 423.840000 ;
      RECT 283.620000 422.760000 326.820000 423.840000 ;
      RECT 238.620000 422.760000 281.820000 423.840000 ;
      RECT 193.620000 422.760000 236.820000 423.840000 ;
      RECT 148.620000 422.760000 191.820000 423.840000 ;
      RECT 103.620000 422.760000 146.820000 423.840000 ;
      RECT 58.620000 422.760000 101.820000 423.840000 ;
      RECT 13.620000 422.760000 56.820000 423.840000 ;
      RECT 7.860000 422.760000 11.820000 423.840000 ;
      RECT 0.000000 422.760000 5.260000 423.840000 ;
      RECT 0.000000 421.900000 548.960000 422.760000 ;
      RECT 0.000000 421.120000 550.160000 421.900000 ;
      RECT 547.900000 420.440000 550.160000 421.120000 ;
      RECT 547.900000 420.040000 548.960000 420.440000 ;
      RECT 506.620000 420.040000 545.300000 421.120000 ;
      RECT 461.620000 420.040000 504.820000 421.120000 ;
      RECT 416.620000 420.040000 459.820000 421.120000 ;
      RECT 371.620000 420.040000 414.820000 421.120000 ;
      RECT 326.620000 420.040000 369.820000 421.120000 ;
      RECT 281.620000 420.040000 324.820000 421.120000 ;
      RECT 236.620000 420.040000 279.820000 421.120000 ;
      RECT 191.620000 420.040000 234.820000 421.120000 ;
      RECT 146.620000 420.040000 189.820000 421.120000 ;
      RECT 101.620000 420.040000 144.820000 421.120000 ;
      RECT 56.620000 420.040000 99.820000 421.120000 ;
      RECT 11.620000 420.040000 54.820000 421.120000 ;
      RECT 4.860000 420.040000 9.655000 421.120000 ;
      RECT 0.000000 420.040000 2.260000 421.120000 ;
      RECT 0.000000 419.460000 548.960000 420.040000 ;
      RECT 0.000000 418.400000 550.160000 419.460000 ;
      RECT 544.900000 418.000000 550.160000 418.400000 ;
      RECT 544.900000 417.320000 548.960000 418.000000 ;
      RECT 508.620000 417.320000 542.300000 418.400000 ;
      RECT 463.620000 417.320000 506.820000 418.400000 ;
      RECT 418.620000 417.320000 461.820000 418.400000 ;
      RECT 373.620000 417.320000 416.820000 418.400000 ;
      RECT 328.620000 417.320000 371.820000 418.400000 ;
      RECT 283.620000 417.320000 326.820000 418.400000 ;
      RECT 238.620000 417.320000 281.820000 418.400000 ;
      RECT 193.620000 417.320000 236.820000 418.400000 ;
      RECT 148.620000 417.320000 191.820000 418.400000 ;
      RECT 103.620000 417.320000 146.820000 418.400000 ;
      RECT 58.620000 417.320000 101.820000 418.400000 ;
      RECT 13.620000 417.320000 56.820000 418.400000 ;
      RECT 7.860000 417.320000 11.820000 418.400000 ;
      RECT 0.000000 417.320000 5.260000 418.400000 ;
      RECT 0.000000 417.020000 548.960000 417.320000 ;
      RECT 0.000000 416.170000 550.160000 417.020000 ;
      RECT 0.000000 415.680000 548.960000 416.170000 ;
      RECT 547.900000 415.190000 548.960000 415.680000 ;
      RECT 547.900000 414.600000 550.160000 415.190000 ;
      RECT 506.620000 414.600000 545.300000 415.680000 ;
      RECT 461.620000 414.600000 504.820000 415.680000 ;
      RECT 416.620000 414.600000 459.820000 415.680000 ;
      RECT 371.620000 414.600000 414.820000 415.680000 ;
      RECT 326.620000 414.600000 369.820000 415.680000 ;
      RECT 281.620000 414.600000 324.820000 415.680000 ;
      RECT 236.620000 414.600000 279.820000 415.680000 ;
      RECT 191.620000 414.600000 234.820000 415.680000 ;
      RECT 146.620000 414.600000 189.820000 415.680000 ;
      RECT 101.620000 414.600000 144.820000 415.680000 ;
      RECT 56.620000 414.600000 99.820000 415.680000 ;
      RECT 11.620000 414.600000 54.820000 415.680000 ;
      RECT 4.860000 414.600000 9.655000 415.680000 ;
      RECT 0.000000 414.600000 2.260000 415.680000 ;
      RECT 0.000000 413.730000 550.160000 414.600000 ;
      RECT 0.000000 412.960000 548.960000 413.730000 ;
      RECT 544.900000 412.750000 548.960000 412.960000 ;
      RECT 544.900000 411.880000 550.160000 412.750000 ;
      RECT 508.620000 411.880000 542.300000 412.960000 ;
      RECT 463.620000 411.880000 506.820000 412.960000 ;
      RECT 418.620000 411.880000 461.820000 412.960000 ;
      RECT 373.620000 411.880000 416.820000 412.960000 ;
      RECT 328.620000 411.880000 371.820000 412.960000 ;
      RECT 283.620000 411.880000 326.820000 412.960000 ;
      RECT 238.620000 411.880000 281.820000 412.960000 ;
      RECT 193.620000 411.880000 236.820000 412.960000 ;
      RECT 148.620000 411.880000 191.820000 412.960000 ;
      RECT 103.620000 411.880000 146.820000 412.960000 ;
      RECT 58.620000 411.880000 101.820000 412.960000 ;
      RECT 13.620000 411.880000 56.820000 412.960000 ;
      RECT 7.860000 411.880000 11.820000 412.960000 ;
      RECT 0.000000 411.880000 5.260000 412.960000 ;
      RECT 0.000000 411.290000 550.160000 411.880000 ;
      RECT 0.000000 410.310000 548.960000 411.290000 ;
      RECT 0.000000 410.240000 550.160000 410.310000 ;
      RECT 547.900000 409.160000 550.160000 410.240000 ;
      RECT 506.620000 409.160000 545.300000 410.240000 ;
      RECT 461.620000 409.160000 504.820000 410.240000 ;
      RECT 416.620000 409.160000 459.820000 410.240000 ;
      RECT 371.620000 409.160000 414.820000 410.240000 ;
      RECT 326.620000 409.160000 369.820000 410.240000 ;
      RECT 281.620000 409.160000 324.820000 410.240000 ;
      RECT 236.620000 409.160000 279.820000 410.240000 ;
      RECT 191.620000 409.160000 234.820000 410.240000 ;
      RECT 146.620000 409.160000 189.820000 410.240000 ;
      RECT 101.620000 409.160000 144.820000 410.240000 ;
      RECT 56.620000 409.160000 99.820000 410.240000 ;
      RECT 11.620000 409.160000 54.820000 410.240000 ;
      RECT 4.860000 409.160000 9.655000 410.240000 ;
      RECT 0.000000 409.160000 2.260000 410.240000 ;
      RECT 0.000000 408.850000 550.160000 409.160000 ;
      RECT 0.000000 407.870000 548.960000 408.850000 ;
      RECT 0.000000 407.520000 550.160000 407.870000 ;
      RECT 544.900000 407.020000 550.160000 407.520000 ;
      RECT 544.900000 406.440000 548.960000 407.020000 ;
      RECT 508.620000 406.440000 542.300000 407.520000 ;
      RECT 463.620000 406.440000 506.820000 407.520000 ;
      RECT 418.620000 406.440000 461.820000 407.520000 ;
      RECT 373.620000 406.440000 416.820000 407.520000 ;
      RECT 328.620000 406.440000 371.820000 407.520000 ;
      RECT 283.620000 406.440000 326.820000 407.520000 ;
      RECT 238.620000 406.440000 281.820000 407.520000 ;
      RECT 193.620000 406.440000 236.820000 407.520000 ;
      RECT 148.620000 406.440000 191.820000 407.520000 ;
      RECT 103.620000 406.440000 146.820000 407.520000 ;
      RECT 58.620000 406.440000 101.820000 407.520000 ;
      RECT 13.620000 406.440000 56.820000 407.520000 ;
      RECT 7.860000 406.440000 11.820000 407.520000 ;
      RECT 0.000000 406.440000 5.260000 407.520000 ;
      RECT 0.000000 406.040000 548.960000 406.440000 ;
      RECT 0.000000 404.800000 550.160000 406.040000 ;
      RECT 547.900000 404.580000 550.160000 404.800000 ;
      RECT 547.900000 403.720000 548.960000 404.580000 ;
      RECT 506.620000 403.720000 545.300000 404.800000 ;
      RECT 461.620000 403.720000 504.820000 404.800000 ;
      RECT 416.620000 403.720000 459.820000 404.800000 ;
      RECT 371.620000 403.720000 414.820000 404.800000 ;
      RECT 326.620000 403.720000 369.820000 404.800000 ;
      RECT 281.620000 403.720000 324.820000 404.800000 ;
      RECT 236.620000 403.720000 279.820000 404.800000 ;
      RECT 191.620000 403.720000 234.820000 404.800000 ;
      RECT 146.620000 403.720000 189.820000 404.800000 ;
      RECT 101.620000 403.720000 144.820000 404.800000 ;
      RECT 56.620000 403.720000 99.820000 404.800000 ;
      RECT 11.620000 403.720000 54.820000 404.800000 ;
      RECT 4.860000 403.720000 9.655000 404.800000 ;
      RECT 0.000000 403.720000 2.260000 404.800000 ;
      RECT 0.000000 403.600000 548.960000 403.720000 ;
      RECT 0.000000 402.140000 550.160000 403.600000 ;
      RECT 0.000000 402.080000 548.960000 402.140000 ;
      RECT 544.900000 401.160000 548.960000 402.080000 ;
      RECT 544.900000 401.000000 550.160000 401.160000 ;
      RECT 508.620000 401.000000 542.300000 402.080000 ;
      RECT 463.620000 401.000000 506.820000 402.080000 ;
      RECT 418.620000 401.000000 461.820000 402.080000 ;
      RECT 373.620000 401.000000 416.820000 402.080000 ;
      RECT 328.620000 401.000000 371.820000 402.080000 ;
      RECT 283.620000 401.000000 326.820000 402.080000 ;
      RECT 238.620000 401.000000 281.820000 402.080000 ;
      RECT 193.620000 401.000000 236.820000 402.080000 ;
      RECT 148.620000 401.000000 191.820000 402.080000 ;
      RECT 103.620000 401.000000 146.820000 402.080000 ;
      RECT 58.620000 401.000000 101.820000 402.080000 ;
      RECT 13.620000 401.000000 56.820000 402.080000 ;
      RECT 7.860000 401.000000 11.820000 402.080000 ;
      RECT 0.000000 401.000000 5.260000 402.080000 ;
      RECT 0.000000 399.700000 550.160000 401.000000 ;
      RECT 0.000000 399.360000 548.960000 399.700000 ;
      RECT 547.900000 398.720000 548.960000 399.360000 ;
      RECT 547.900000 398.280000 550.160000 398.720000 ;
      RECT 506.620000 398.280000 545.300000 399.360000 ;
      RECT 461.620000 398.280000 504.820000 399.360000 ;
      RECT 416.620000 398.280000 459.820000 399.360000 ;
      RECT 371.620000 398.280000 414.820000 399.360000 ;
      RECT 326.620000 398.280000 369.820000 399.360000 ;
      RECT 281.620000 398.280000 324.820000 399.360000 ;
      RECT 236.620000 398.280000 279.820000 399.360000 ;
      RECT 191.620000 398.280000 234.820000 399.360000 ;
      RECT 146.620000 398.280000 189.820000 399.360000 ;
      RECT 101.620000 398.280000 144.820000 399.360000 ;
      RECT 56.620000 398.280000 99.820000 399.360000 ;
      RECT 11.620000 398.280000 54.820000 399.360000 ;
      RECT 4.860000 398.280000 9.655000 399.360000 ;
      RECT 0.000000 398.280000 2.260000 399.360000 ;
      RECT 0.000000 397.870000 550.160000 398.280000 ;
      RECT 0.000000 396.890000 548.960000 397.870000 ;
      RECT 0.000000 396.640000 550.160000 396.890000 ;
      RECT 544.900000 395.560000 550.160000 396.640000 ;
      RECT 508.620000 395.560000 542.300000 396.640000 ;
      RECT 463.620000 395.560000 506.820000 396.640000 ;
      RECT 418.620000 395.560000 461.820000 396.640000 ;
      RECT 373.620000 395.560000 416.820000 396.640000 ;
      RECT 328.620000 395.560000 371.820000 396.640000 ;
      RECT 283.620000 395.560000 326.820000 396.640000 ;
      RECT 238.620000 395.560000 281.820000 396.640000 ;
      RECT 193.620000 395.560000 236.820000 396.640000 ;
      RECT 148.620000 395.560000 191.820000 396.640000 ;
      RECT 103.620000 395.560000 146.820000 396.640000 ;
      RECT 58.620000 395.560000 101.820000 396.640000 ;
      RECT 13.620000 395.560000 56.820000 396.640000 ;
      RECT 7.860000 395.560000 11.820000 396.640000 ;
      RECT 0.000000 395.560000 5.260000 396.640000 ;
      RECT 0.000000 395.430000 550.160000 395.560000 ;
      RECT 0.000000 394.450000 548.960000 395.430000 ;
      RECT 0.000000 393.920000 550.160000 394.450000 ;
      RECT 547.900000 392.990000 550.160000 393.920000 ;
      RECT 547.900000 392.840000 548.960000 392.990000 ;
      RECT 506.620000 392.840000 545.300000 393.920000 ;
      RECT 461.620000 392.840000 504.820000 393.920000 ;
      RECT 416.620000 392.840000 459.820000 393.920000 ;
      RECT 371.620000 392.840000 414.820000 393.920000 ;
      RECT 326.620000 392.840000 369.820000 393.920000 ;
      RECT 281.620000 392.840000 324.820000 393.920000 ;
      RECT 236.620000 392.840000 279.820000 393.920000 ;
      RECT 191.620000 392.840000 234.820000 393.920000 ;
      RECT 146.620000 392.840000 189.820000 393.920000 ;
      RECT 101.620000 392.840000 144.820000 393.920000 ;
      RECT 56.620000 392.840000 99.820000 393.920000 ;
      RECT 11.620000 392.840000 54.820000 393.920000 ;
      RECT 4.860000 392.840000 9.655000 393.920000 ;
      RECT 0.000000 392.840000 2.260000 393.920000 ;
      RECT 0.000000 392.010000 548.960000 392.840000 ;
      RECT 0.000000 391.200000 550.160000 392.010000 ;
      RECT 544.900000 390.550000 550.160000 391.200000 ;
      RECT 544.900000 390.120000 548.960000 390.550000 ;
      RECT 508.620000 390.120000 542.300000 391.200000 ;
      RECT 463.620000 390.120000 506.820000 391.200000 ;
      RECT 418.620000 390.120000 461.820000 391.200000 ;
      RECT 373.620000 390.120000 416.820000 391.200000 ;
      RECT 328.620000 390.120000 371.820000 391.200000 ;
      RECT 283.620000 390.120000 326.820000 391.200000 ;
      RECT 238.620000 390.120000 281.820000 391.200000 ;
      RECT 193.620000 390.120000 236.820000 391.200000 ;
      RECT 148.620000 390.120000 191.820000 391.200000 ;
      RECT 103.620000 390.120000 146.820000 391.200000 ;
      RECT 58.620000 390.120000 101.820000 391.200000 ;
      RECT 13.620000 390.120000 56.820000 391.200000 ;
      RECT 7.860000 390.120000 11.820000 391.200000 ;
      RECT 0.000000 390.120000 5.260000 391.200000 ;
      RECT 0.000000 389.570000 548.960000 390.120000 ;
      RECT 0.000000 388.480000 550.160000 389.570000 ;
      RECT 547.900000 388.110000 550.160000 388.480000 ;
      RECT 547.900000 387.400000 548.960000 388.110000 ;
      RECT 506.620000 387.400000 545.300000 388.480000 ;
      RECT 461.620000 387.400000 504.820000 388.480000 ;
      RECT 416.620000 387.400000 459.820000 388.480000 ;
      RECT 371.620000 387.400000 414.820000 388.480000 ;
      RECT 326.620000 387.400000 369.820000 388.480000 ;
      RECT 281.620000 387.400000 324.820000 388.480000 ;
      RECT 236.620000 387.400000 279.820000 388.480000 ;
      RECT 191.620000 387.400000 234.820000 388.480000 ;
      RECT 146.620000 387.400000 189.820000 388.480000 ;
      RECT 101.620000 387.400000 144.820000 388.480000 ;
      RECT 56.620000 387.400000 99.820000 388.480000 ;
      RECT 11.620000 387.400000 54.820000 388.480000 ;
      RECT 4.860000 387.400000 9.655000 388.480000 ;
      RECT 0.000000 387.400000 2.260000 388.480000 ;
      RECT 0.000000 387.130000 548.960000 387.400000 ;
      RECT 0.000000 386.280000 550.160000 387.130000 ;
      RECT 0.000000 385.760000 548.960000 386.280000 ;
      RECT 544.900000 385.300000 548.960000 385.760000 ;
      RECT 544.900000 384.680000 550.160000 385.300000 ;
      RECT 508.620000 384.680000 542.300000 385.760000 ;
      RECT 463.620000 384.680000 506.820000 385.760000 ;
      RECT 418.620000 384.680000 461.820000 385.760000 ;
      RECT 373.620000 384.680000 416.820000 385.760000 ;
      RECT 328.620000 384.680000 371.820000 385.760000 ;
      RECT 283.620000 384.680000 326.820000 385.760000 ;
      RECT 238.620000 384.680000 281.820000 385.760000 ;
      RECT 193.620000 384.680000 236.820000 385.760000 ;
      RECT 148.620000 384.680000 191.820000 385.760000 ;
      RECT 103.620000 384.680000 146.820000 385.760000 ;
      RECT 58.620000 384.680000 101.820000 385.760000 ;
      RECT 13.620000 384.680000 56.820000 385.760000 ;
      RECT 7.860000 384.680000 11.820000 385.760000 ;
      RECT 0.000000 384.680000 5.260000 385.760000 ;
      RECT 0.000000 383.840000 550.160000 384.680000 ;
      RECT 0.000000 383.040000 548.960000 383.840000 ;
      RECT 547.900000 382.860000 548.960000 383.040000 ;
      RECT 547.900000 381.960000 550.160000 382.860000 ;
      RECT 506.620000 381.960000 545.300000 383.040000 ;
      RECT 461.620000 381.960000 504.820000 383.040000 ;
      RECT 416.620000 381.960000 459.820000 383.040000 ;
      RECT 371.620000 381.960000 414.820000 383.040000 ;
      RECT 326.620000 381.960000 369.820000 383.040000 ;
      RECT 281.620000 381.960000 324.820000 383.040000 ;
      RECT 236.620000 381.960000 279.820000 383.040000 ;
      RECT 191.620000 381.960000 234.820000 383.040000 ;
      RECT 146.620000 381.960000 189.820000 383.040000 ;
      RECT 101.620000 381.960000 144.820000 383.040000 ;
      RECT 56.620000 381.960000 99.820000 383.040000 ;
      RECT 11.620000 381.960000 54.820000 383.040000 ;
      RECT 4.860000 381.960000 9.655000 383.040000 ;
      RECT 0.000000 381.960000 2.260000 383.040000 ;
      RECT 0.000000 381.400000 550.160000 381.960000 ;
      RECT 0.000000 380.420000 548.960000 381.400000 ;
      RECT 0.000000 380.320000 550.160000 380.420000 ;
      RECT 544.900000 379.240000 550.160000 380.320000 ;
      RECT 508.620000 379.240000 542.300000 380.320000 ;
      RECT 463.620000 379.240000 506.820000 380.320000 ;
      RECT 418.620000 379.240000 461.820000 380.320000 ;
      RECT 373.620000 379.240000 416.820000 380.320000 ;
      RECT 328.620000 379.240000 371.820000 380.320000 ;
      RECT 283.620000 379.240000 326.820000 380.320000 ;
      RECT 238.620000 379.240000 281.820000 380.320000 ;
      RECT 193.620000 379.240000 236.820000 380.320000 ;
      RECT 148.620000 379.240000 191.820000 380.320000 ;
      RECT 103.620000 379.240000 146.820000 380.320000 ;
      RECT 58.620000 379.240000 101.820000 380.320000 ;
      RECT 13.620000 379.240000 56.820000 380.320000 ;
      RECT 7.860000 379.240000 11.820000 380.320000 ;
      RECT 0.000000 379.240000 5.260000 380.320000 ;
      RECT 0.000000 378.960000 550.160000 379.240000 ;
      RECT 0.000000 377.980000 548.960000 378.960000 ;
      RECT 0.000000 377.600000 550.160000 377.980000 ;
      RECT 547.900000 377.130000 550.160000 377.600000 ;
      RECT 547.900000 376.520000 548.960000 377.130000 ;
      RECT 506.620000 376.520000 545.300000 377.600000 ;
      RECT 461.620000 376.520000 504.820000 377.600000 ;
      RECT 416.620000 376.520000 459.820000 377.600000 ;
      RECT 371.620000 376.520000 414.820000 377.600000 ;
      RECT 326.620000 376.520000 369.820000 377.600000 ;
      RECT 281.620000 376.520000 324.820000 377.600000 ;
      RECT 236.620000 376.520000 279.820000 377.600000 ;
      RECT 191.620000 376.520000 234.820000 377.600000 ;
      RECT 146.620000 376.520000 189.820000 377.600000 ;
      RECT 101.620000 376.520000 144.820000 377.600000 ;
      RECT 56.620000 376.520000 99.820000 377.600000 ;
      RECT 11.620000 376.520000 54.820000 377.600000 ;
      RECT 4.860000 376.520000 9.655000 377.600000 ;
      RECT 0.000000 376.520000 2.260000 377.600000 ;
      RECT 0.000000 376.150000 548.960000 376.520000 ;
      RECT 0.000000 374.880000 550.160000 376.150000 ;
      RECT 544.900000 374.690000 550.160000 374.880000 ;
      RECT 544.900000 373.800000 548.960000 374.690000 ;
      RECT 508.620000 373.800000 542.300000 374.880000 ;
      RECT 463.620000 373.800000 506.820000 374.880000 ;
      RECT 418.620000 373.800000 461.820000 374.880000 ;
      RECT 373.620000 373.800000 416.820000 374.880000 ;
      RECT 328.620000 373.800000 371.820000 374.880000 ;
      RECT 283.620000 373.800000 326.820000 374.880000 ;
      RECT 238.620000 373.800000 281.820000 374.880000 ;
      RECT 193.620000 373.800000 236.820000 374.880000 ;
      RECT 148.620000 373.800000 191.820000 374.880000 ;
      RECT 103.620000 373.800000 146.820000 374.880000 ;
      RECT 58.620000 373.800000 101.820000 374.880000 ;
      RECT 13.620000 373.800000 56.820000 374.880000 ;
      RECT 7.860000 373.800000 11.820000 374.880000 ;
      RECT 0.000000 373.800000 5.260000 374.880000 ;
      RECT 0.000000 373.710000 548.960000 373.800000 ;
      RECT 0.000000 372.250000 550.160000 373.710000 ;
      RECT 0.000000 372.160000 548.960000 372.250000 ;
      RECT 547.900000 371.270000 548.960000 372.160000 ;
      RECT 547.900000 371.080000 550.160000 371.270000 ;
      RECT 506.620000 371.080000 545.300000 372.160000 ;
      RECT 461.620000 371.080000 504.820000 372.160000 ;
      RECT 416.620000 371.080000 459.820000 372.160000 ;
      RECT 371.620000 371.080000 414.820000 372.160000 ;
      RECT 326.620000 371.080000 369.820000 372.160000 ;
      RECT 281.620000 371.080000 324.820000 372.160000 ;
      RECT 236.620000 371.080000 279.820000 372.160000 ;
      RECT 191.620000 371.080000 234.820000 372.160000 ;
      RECT 146.620000 371.080000 189.820000 372.160000 ;
      RECT 101.620000 371.080000 144.820000 372.160000 ;
      RECT 56.620000 371.080000 99.820000 372.160000 ;
      RECT 11.620000 371.080000 54.820000 372.160000 ;
      RECT 4.860000 371.080000 9.655000 372.160000 ;
      RECT 0.000000 371.080000 2.260000 372.160000 ;
      RECT 0.000000 369.810000 550.160000 371.080000 ;
      RECT 0.000000 369.440000 548.960000 369.810000 ;
      RECT 544.900000 368.830000 548.960000 369.440000 ;
      RECT 544.900000 368.360000 550.160000 368.830000 ;
      RECT 508.620000 368.360000 542.300000 369.440000 ;
      RECT 463.620000 368.360000 506.820000 369.440000 ;
      RECT 418.620000 368.360000 461.820000 369.440000 ;
      RECT 373.620000 368.360000 416.820000 369.440000 ;
      RECT 328.620000 368.360000 371.820000 369.440000 ;
      RECT 283.620000 368.360000 326.820000 369.440000 ;
      RECT 238.620000 368.360000 281.820000 369.440000 ;
      RECT 193.620000 368.360000 236.820000 369.440000 ;
      RECT 148.620000 368.360000 191.820000 369.440000 ;
      RECT 103.620000 368.360000 146.820000 369.440000 ;
      RECT 58.620000 368.360000 101.820000 369.440000 ;
      RECT 13.620000 368.360000 56.820000 369.440000 ;
      RECT 7.860000 368.360000 11.820000 369.440000 ;
      RECT 0.000000 368.360000 5.260000 369.440000 ;
      RECT 0.000000 367.980000 550.160000 368.360000 ;
      RECT 0.000000 367.000000 548.960000 367.980000 ;
      RECT 0.000000 366.720000 550.160000 367.000000 ;
      RECT 547.900000 365.640000 550.160000 366.720000 ;
      RECT 506.620000 365.640000 545.300000 366.720000 ;
      RECT 461.620000 365.640000 504.820000 366.720000 ;
      RECT 416.620000 365.640000 459.820000 366.720000 ;
      RECT 371.620000 365.640000 414.820000 366.720000 ;
      RECT 326.620000 365.640000 369.820000 366.720000 ;
      RECT 281.620000 365.640000 324.820000 366.720000 ;
      RECT 236.620000 365.640000 279.820000 366.720000 ;
      RECT 191.620000 365.640000 234.820000 366.720000 ;
      RECT 146.620000 365.640000 189.820000 366.720000 ;
      RECT 101.620000 365.640000 144.820000 366.720000 ;
      RECT 56.620000 365.640000 99.820000 366.720000 ;
      RECT 11.620000 365.640000 54.820000 366.720000 ;
      RECT 4.860000 365.640000 9.655000 366.720000 ;
      RECT 0.000000 365.640000 2.260000 366.720000 ;
      RECT 0.000000 365.540000 550.160000 365.640000 ;
      RECT 0.000000 364.560000 548.960000 365.540000 ;
      RECT 0.000000 364.000000 550.160000 364.560000 ;
      RECT 544.900000 363.100000 550.160000 364.000000 ;
      RECT 544.900000 362.920000 548.960000 363.100000 ;
      RECT 508.620000 362.920000 542.300000 364.000000 ;
      RECT 463.620000 362.920000 506.820000 364.000000 ;
      RECT 418.620000 362.920000 461.820000 364.000000 ;
      RECT 373.620000 362.920000 416.820000 364.000000 ;
      RECT 328.620000 362.920000 371.820000 364.000000 ;
      RECT 283.620000 362.920000 326.820000 364.000000 ;
      RECT 238.620000 362.920000 281.820000 364.000000 ;
      RECT 193.620000 362.920000 236.820000 364.000000 ;
      RECT 148.620000 362.920000 191.820000 364.000000 ;
      RECT 103.620000 362.920000 146.820000 364.000000 ;
      RECT 58.620000 362.920000 101.820000 364.000000 ;
      RECT 13.620000 362.920000 56.820000 364.000000 ;
      RECT 7.860000 362.920000 11.820000 364.000000 ;
      RECT 0.000000 362.920000 5.260000 364.000000 ;
      RECT 0.000000 362.120000 548.960000 362.920000 ;
      RECT 0.000000 361.280000 550.160000 362.120000 ;
      RECT 547.900000 360.660000 550.160000 361.280000 ;
      RECT 547.900000 360.200000 548.960000 360.660000 ;
      RECT 506.620000 360.200000 545.300000 361.280000 ;
      RECT 461.620000 360.200000 504.820000 361.280000 ;
      RECT 416.620000 360.200000 459.820000 361.280000 ;
      RECT 371.620000 360.200000 414.820000 361.280000 ;
      RECT 326.620000 360.200000 369.820000 361.280000 ;
      RECT 281.620000 360.200000 324.820000 361.280000 ;
      RECT 236.620000 360.200000 279.820000 361.280000 ;
      RECT 191.620000 360.200000 234.820000 361.280000 ;
      RECT 146.620000 360.200000 189.820000 361.280000 ;
      RECT 101.620000 360.200000 144.820000 361.280000 ;
      RECT 56.620000 360.200000 99.820000 361.280000 ;
      RECT 11.620000 360.200000 54.820000 361.280000 ;
      RECT 4.860000 360.200000 9.655000 361.280000 ;
      RECT 0.000000 360.200000 2.260000 361.280000 ;
      RECT 0.000000 359.680000 548.960000 360.200000 ;
      RECT 0.000000 358.830000 550.160000 359.680000 ;
      RECT 0.000000 358.560000 548.960000 358.830000 ;
      RECT 544.900000 357.850000 548.960000 358.560000 ;
      RECT 544.900000 357.480000 550.160000 357.850000 ;
      RECT 508.620000 357.480000 542.300000 358.560000 ;
      RECT 463.620000 357.480000 506.820000 358.560000 ;
      RECT 418.620000 357.480000 461.820000 358.560000 ;
      RECT 373.620000 357.480000 416.820000 358.560000 ;
      RECT 328.620000 357.480000 371.820000 358.560000 ;
      RECT 283.620000 357.480000 326.820000 358.560000 ;
      RECT 238.620000 357.480000 281.820000 358.560000 ;
      RECT 193.620000 357.480000 236.820000 358.560000 ;
      RECT 148.620000 357.480000 191.820000 358.560000 ;
      RECT 103.620000 357.480000 146.820000 358.560000 ;
      RECT 58.620000 357.480000 101.820000 358.560000 ;
      RECT 13.620000 357.480000 56.820000 358.560000 ;
      RECT 7.860000 357.480000 11.820000 358.560000 ;
      RECT 0.000000 357.480000 5.260000 358.560000 ;
      RECT 0.000000 356.390000 550.160000 357.480000 ;
      RECT 0.000000 355.840000 548.960000 356.390000 ;
      RECT 547.900000 355.410000 548.960000 355.840000 ;
      RECT 547.900000 354.760000 550.160000 355.410000 ;
      RECT 506.620000 354.760000 545.300000 355.840000 ;
      RECT 461.620000 354.760000 504.820000 355.840000 ;
      RECT 416.620000 354.760000 459.820000 355.840000 ;
      RECT 371.620000 354.760000 414.820000 355.840000 ;
      RECT 326.620000 354.760000 369.820000 355.840000 ;
      RECT 281.620000 354.760000 324.820000 355.840000 ;
      RECT 236.620000 354.760000 279.820000 355.840000 ;
      RECT 191.620000 354.760000 234.820000 355.840000 ;
      RECT 146.620000 354.760000 189.820000 355.840000 ;
      RECT 101.620000 354.760000 144.820000 355.840000 ;
      RECT 56.620000 354.760000 99.820000 355.840000 ;
      RECT 11.620000 354.760000 54.820000 355.840000 ;
      RECT 4.860000 354.760000 9.655000 355.840000 ;
      RECT 0.000000 354.760000 2.260000 355.840000 ;
      RECT 0.000000 353.950000 550.160000 354.760000 ;
      RECT 0.000000 353.120000 548.960000 353.950000 ;
      RECT 544.900000 352.970000 548.960000 353.120000 ;
      RECT 544.900000 352.040000 550.160000 352.970000 ;
      RECT 508.620000 352.040000 542.300000 353.120000 ;
      RECT 463.620000 352.040000 506.820000 353.120000 ;
      RECT 418.620000 352.040000 461.820000 353.120000 ;
      RECT 373.620000 352.040000 416.820000 353.120000 ;
      RECT 328.620000 352.040000 371.820000 353.120000 ;
      RECT 283.620000 352.040000 326.820000 353.120000 ;
      RECT 238.620000 352.040000 281.820000 353.120000 ;
      RECT 193.620000 352.040000 236.820000 353.120000 ;
      RECT 148.620000 352.040000 191.820000 353.120000 ;
      RECT 103.620000 352.040000 146.820000 353.120000 ;
      RECT 58.620000 352.040000 101.820000 353.120000 ;
      RECT 13.620000 352.040000 56.820000 353.120000 ;
      RECT 7.860000 352.040000 11.820000 353.120000 ;
      RECT 0.000000 352.040000 5.260000 353.120000 ;
      RECT 0.000000 351.510000 550.160000 352.040000 ;
      RECT 0.000000 350.530000 548.960000 351.510000 ;
      RECT 0.000000 350.400000 550.160000 350.530000 ;
      RECT 547.900000 349.680000 550.160000 350.400000 ;
      RECT 547.900000 349.320000 548.960000 349.680000 ;
      RECT 506.620000 349.320000 545.300000 350.400000 ;
      RECT 461.620000 349.320000 504.820000 350.400000 ;
      RECT 416.620000 349.320000 459.820000 350.400000 ;
      RECT 371.620000 349.320000 414.820000 350.400000 ;
      RECT 326.620000 349.320000 369.820000 350.400000 ;
      RECT 281.620000 349.320000 324.820000 350.400000 ;
      RECT 236.620000 349.320000 279.820000 350.400000 ;
      RECT 191.620000 349.320000 234.820000 350.400000 ;
      RECT 146.620000 349.320000 189.820000 350.400000 ;
      RECT 101.620000 349.320000 144.820000 350.400000 ;
      RECT 56.620000 349.320000 99.820000 350.400000 ;
      RECT 11.620000 349.320000 54.820000 350.400000 ;
      RECT 4.860000 349.320000 9.655000 350.400000 ;
      RECT 0.000000 349.320000 2.260000 350.400000 ;
      RECT 0.000000 348.700000 548.960000 349.320000 ;
      RECT 0.000000 347.680000 550.160000 348.700000 ;
      RECT 544.900000 347.240000 550.160000 347.680000 ;
      RECT 544.900000 346.600000 548.960000 347.240000 ;
      RECT 508.620000 346.600000 542.300000 347.680000 ;
      RECT 463.620000 346.600000 506.820000 347.680000 ;
      RECT 418.620000 346.600000 461.820000 347.680000 ;
      RECT 373.620000 346.600000 416.820000 347.680000 ;
      RECT 328.620000 346.600000 371.820000 347.680000 ;
      RECT 283.620000 346.600000 326.820000 347.680000 ;
      RECT 238.620000 346.600000 281.820000 347.680000 ;
      RECT 193.620000 346.600000 236.820000 347.680000 ;
      RECT 148.620000 346.600000 191.820000 347.680000 ;
      RECT 103.620000 346.600000 146.820000 347.680000 ;
      RECT 58.620000 346.600000 101.820000 347.680000 ;
      RECT 13.620000 346.600000 56.820000 347.680000 ;
      RECT 7.860000 346.600000 11.820000 347.680000 ;
      RECT 0.000000 346.600000 5.260000 347.680000 ;
      RECT 0.000000 346.260000 548.960000 346.600000 ;
      RECT 0.000000 344.960000 550.160000 346.260000 ;
      RECT 547.900000 344.800000 550.160000 344.960000 ;
      RECT 547.900000 343.880000 548.960000 344.800000 ;
      RECT 506.620000 343.880000 545.300000 344.960000 ;
      RECT 461.620000 343.880000 504.820000 344.960000 ;
      RECT 416.620000 343.880000 459.820000 344.960000 ;
      RECT 371.620000 343.880000 414.820000 344.960000 ;
      RECT 326.620000 343.880000 369.820000 344.960000 ;
      RECT 281.620000 343.880000 324.820000 344.960000 ;
      RECT 236.620000 343.880000 279.820000 344.960000 ;
      RECT 191.620000 343.880000 234.820000 344.960000 ;
      RECT 146.620000 343.880000 189.820000 344.960000 ;
      RECT 101.620000 343.880000 144.820000 344.960000 ;
      RECT 56.620000 343.880000 99.820000 344.960000 ;
      RECT 11.620000 343.880000 54.820000 344.960000 ;
      RECT 4.860000 343.880000 9.655000 344.960000 ;
      RECT 0.000000 343.880000 2.260000 344.960000 ;
      RECT 0.000000 343.820000 548.960000 343.880000 ;
      RECT 0.000000 342.360000 550.160000 343.820000 ;
      RECT 0.000000 342.240000 548.960000 342.360000 ;
      RECT 544.900000 341.380000 548.960000 342.240000 ;
      RECT 544.900000 341.160000 550.160000 341.380000 ;
      RECT 508.620000 341.160000 542.300000 342.240000 ;
      RECT 463.620000 341.160000 506.820000 342.240000 ;
      RECT 418.620000 341.160000 461.820000 342.240000 ;
      RECT 373.620000 341.160000 416.820000 342.240000 ;
      RECT 328.620000 341.160000 371.820000 342.240000 ;
      RECT 283.620000 341.160000 326.820000 342.240000 ;
      RECT 238.620000 341.160000 281.820000 342.240000 ;
      RECT 193.620000 341.160000 236.820000 342.240000 ;
      RECT 148.620000 341.160000 191.820000 342.240000 ;
      RECT 103.620000 341.160000 146.820000 342.240000 ;
      RECT 58.620000 341.160000 101.820000 342.240000 ;
      RECT 13.620000 341.160000 56.820000 342.240000 ;
      RECT 7.860000 341.160000 11.820000 342.240000 ;
      RECT 0.000000 341.160000 5.260000 342.240000 ;
      RECT 0.000000 340.530000 550.160000 341.160000 ;
      RECT 0.000000 339.550000 548.960000 340.530000 ;
      RECT 0.000000 339.520000 550.160000 339.550000 ;
      RECT 547.900000 338.440000 550.160000 339.520000 ;
      RECT 506.620000 338.440000 545.300000 339.520000 ;
      RECT 461.620000 338.440000 504.820000 339.520000 ;
      RECT 416.620000 338.440000 459.820000 339.520000 ;
      RECT 371.620000 338.440000 414.820000 339.520000 ;
      RECT 326.620000 338.440000 369.820000 339.520000 ;
      RECT 281.620000 338.440000 324.820000 339.520000 ;
      RECT 236.620000 338.440000 279.820000 339.520000 ;
      RECT 191.620000 338.440000 234.820000 339.520000 ;
      RECT 146.620000 338.440000 189.820000 339.520000 ;
      RECT 101.620000 338.440000 144.820000 339.520000 ;
      RECT 56.620000 338.440000 99.820000 339.520000 ;
      RECT 11.620000 338.440000 54.820000 339.520000 ;
      RECT 4.860000 338.440000 9.655000 339.520000 ;
      RECT 0.000000 338.440000 2.260000 339.520000 ;
      RECT 0.000000 338.090000 550.160000 338.440000 ;
      RECT 0.000000 337.110000 548.960000 338.090000 ;
      RECT 0.000000 336.800000 550.160000 337.110000 ;
      RECT 544.900000 335.720000 550.160000 336.800000 ;
      RECT 508.620000 335.720000 542.300000 336.800000 ;
      RECT 463.620000 335.720000 506.820000 336.800000 ;
      RECT 418.620000 335.720000 461.820000 336.800000 ;
      RECT 373.620000 335.720000 416.820000 336.800000 ;
      RECT 328.620000 335.720000 371.820000 336.800000 ;
      RECT 283.620000 335.720000 326.820000 336.800000 ;
      RECT 238.620000 335.720000 281.820000 336.800000 ;
      RECT 193.620000 335.720000 236.820000 336.800000 ;
      RECT 148.620000 335.720000 191.820000 336.800000 ;
      RECT 103.620000 335.720000 146.820000 336.800000 ;
      RECT 58.620000 335.720000 101.820000 336.800000 ;
      RECT 13.620000 335.720000 56.820000 336.800000 ;
      RECT 7.860000 335.720000 11.820000 336.800000 ;
      RECT 0.000000 335.720000 5.260000 336.800000 ;
      RECT 0.000000 335.650000 550.160000 335.720000 ;
      RECT 0.000000 334.670000 548.960000 335.650000 ;
      RECT 0.000000 334.080000 550.160000 334.670000 ;
      RECT 547.900000 333.210000 550.160000 334.080000 ;
      RECT 547.900000 333.000000 548.960000 333.210000 ;
      RECT 506.620000 333.000000 545.300000 334.080000 ;
      RECT 461.620000 333.000000 504.820000 334.080000 ;
      RECT 416.620000 333.000000 459.820000 334.080000 ;
      RECT 371.620000 333.000000 414.820000 334.080000 ;
      RECT 326.620000 333.000000 369.820000 334.080000 ;
      RECT 281.620000 333.000000 324.820000 334.080000 ;
      RECT 236.620000 333.000000 279.820000 334.080000 ;
      RECT 191.620000 333.000000 234.820000 334.080000 ;
      RECT 146.620000 333.000000 189.820000 334.080000 ;
      RECT 101.620000 333.000000 144.820000 334.080000 ;
      RECT 56.620000 333.000000 99.820000 334.080000 ;
      RECT 11.620000 333.000000 54.820000 334.080000 ;
      RECT 4.860000 333.000000 9.655000 334.080000 ;
      RECT 0.000000 333.000000 2.260000 334.080000 ;
      RECT 0.000000 332.230000 548.960000 333.000000 ;
      RECT 0.000000 331.380000 550.160000 332.230000 ;
      RECT 0.000000 331.360000 548.960000 331.380000 ;
      RECT 544.900000 330.400000 548.960000 331.360000 ;
      RECT 544.900000 330.280000 550.160000 330.400000 ;
      RECT 508.620000 330.280000 542.300000 331.360000 ;
      RECT 463.620000 330.280000 506.820000 331.360000 ;
      RECT 418.620000 330.280000 461.820000 331.360000 ;
      RECT 373.620000 330.280000 416.820000 331.360000 ;
      RECT 328.620000 330.280000 371.820000 331.360000 ;
      RECT 283.620000 330.280000 326.820000 331.360000 ;
      RECT 238.620000 330.280000 281.820000 331.360000 ;
      RECT 193.620000 330.280000 236.820000 331.360000 ;
      RECT 148.620000 330.280000 191.820000 331.360000 ;
      RECT 103.620000 330.280000 146.820000 331.360000 ;
      RECT 58.620000 330.280000 101.820000 331.360000 ;
      RECT 13.620000 330.280000 56.820000 331.360000 ;
      RECT 7.860000 330.280000 11.820000 331.360000 ;
      RECT 0.000000 330.280000 5.260000 331.360000 ;
      RECT 0.000000 328.940000 550.160000 330.280000 ;
      RECT 0.000000 328.640000 548.960000 328.940000 ;
      RECT 547.900000 327.960000 548.960000 328.640000 ;
      RECT 547.900000 327.560000 550.160000 327.960000 ;
      RECT 506.620000 327.560000 545.300000 328.640000 ;
      RECT 461.620000 327.560000 504.820000 328.640000 ;
      RECT 416.620000 327.560000 459.820000 328.640000 ;
      RECT 371.620000 327.560000 414.820000 328.640000 ;
      RECT 326.620000 327.560000 369.820000 328.640000 ;
      RECT 281.620000 327.560000 324.820000 328.640000 ;
      RECT 236.620000 327.560000 279.820000 328.640000 ;
      RECT 191.620000 327.560000 234.820000 328.640000 ;
      RECT 146.620000 327.560000 189.820000 328.640000 ;
      RECT 101.620000 327.560000 144.820000 328.640000 ;
      RECT 56.620000 327.560000 99.820000 328.640000 ;
      RECT 11.620000 327.560000 54.820000 328.640000 ;
      RECT 4.860000 327.560000 9.655000 328.640000 ;
      RECT 0.000000 327.560000 2.260000 328.640000 ;
      RECT 0.000000 326.500000 550.160000 327.560000 ;
      RECT 0.000000 325.920000 548.960000 326.500000 ;
      RECT 544.900000 325.520000 548.960000 325.920000 ;
      RECT 544.900000 324.840000 550.160000 325.520000 ;
      RECT 508.620000 324.840000 542.300000 325.920000 ;
      RECT 463.620000 324.840000 506.820000 325.920000 ;
      RECT 418.620000 324.840000 461.820000 325.920000 ;
      RECT 373.620000 324.840000 416.820000 325.920000 ;
      RECT 328.620000 324.840000 371.820000 325.920000 ;
      RECT 283.620000 324.840000 326.820000 325.920000 ;
      RECT 238.620000 324.840000 281.820000 325.920000 ;
      RECT 193.620000 324.840000 236.820000 325.920000 ;
      RECT 148.620000 324.840000 191.820000 325.920000 ;
      RECT 103.620000 324.840000 146.820000 325.920000 ;
      RECT 58.620000 324.840000 101.820000 325.920000 ;
      RECT 13.620000 324.840000 56.820000 325.920000 ;
      RECT 7.860000 324.840000 11.820000 325.920000 ;
      RECT 0.000000 324.840000 5.260000 325.920000 ;
      RECT 0.000000 324.060000 550.160000 324.840000 ;
      RECT 0.000000 323.200000 548.960000 324.060000 ;
      RECT 547.900000 323.080000 548.960000 323.200000 ;
      RECT 547.900000 322.230000 550.160000 323.080000 ;
      RECT 547.900000 322.120000 548.960000 322.230000 ;
      RECT 506.620000 322.120000 545.300000 323.200000 ;
      RECT 461.620000 322.120000 504.820000 323.200000 ;
      RECT 416.620000 322.120000 459.820000 323.200000 ;
      RECT 371.620000 322.120000 414.820000 323.200000 ;
      RECT 326.620000 322.120000 369.820000 323.200000 ;
      RECT 281.620000 322.120000 324.820000 323.200000 ;
      RECT 236.620000 322.120000 279.820000 323.200000 ;
      RECT 191.620000 322.120000 234.820000 323.200000 ;
      RECT 146.620000 322.120000 189.820000 323.200000 ;
      RECT 101.620000 322.120000 144.820000 323.200000 ;
      RECT 56.620000 322.120000 99.820000 323.200000 ;
      RECT 11.620000 322.120000 54.820000 323.200000 ;
      RECT 4.860000 322.120000 9.655000 323.200000 ;
      RECT 0.000000 322.120000 2.260000 323.200000 ;
      RECT 0.000000 321.250000 548.960000 322.120000 ;
      RECT 0.000000 320.480000 550.160000 321.250000 ;
      RECT 544.900000 319.790000 550.160000 320.480000 ;
      RECT 544.900000 319.400000 548.960000 319.790000 ;
      RECT 508.620000 319.400000 542.300000 320.480000 ;
      RECT 463.620000 319.400000 506.820000 320.480000 ;
      RECT 418.620000 319.400000 461.820000 320.480000 ;
      RECT 373.620000 319.400000 416.820000 320.480000 ;
      RECT 328.620000 319.400000 371.820000 320.480000 ;
      RECT 283.620000 319.400000 326.820000 320.480000 ;
      RECT 238.620000 319.400000 281.820000 320.480000 ;
      RECT 193.620000 319.400000 236.820000 320.480000 ;
      RECT 148.620000 319.400000 191.820000 320.480000 ;
      RECT 103.620000 319.400000 146.820000 320.480000 ;
      RECT 58.620000 319.400000 101.820000 320.480000 ;
      RECT 13.620000 319.400000 56.820000 320.480000 ;
      RECT 7.860000 319.400000 11.820000 320.480000 ;
      RECT 0.000000 319.400000 5.260000 320.480000 ;
      RECT 0.000000 318.810000 548.960000 319.400000 ;
      RECT 0.000000 317.760000 550.160000 318.810000 ;
      RECT 547.900000 317.350000 550.160000 317.760000 ;
      RECT 547.900000 316.680000 548.960000 317.350000 ;
      RECT 506.620000 316.680000 545.300000 317.760000 ;
      RECT 461.620000 316.680000 504.820000 317.760000 ;
      RECT 416.620000 316.680000 459.820000 317.760000 ;
      RECT 371.620000 316.680000 414.820000 317.760000 ;
      RECT 326.620000 316.680000 369.820000 317.760000 ;
      RECT 281.620000 316.680000 324.820000 317.760000 ;
      RECT 236.620000 316.680000 279.820000 317.760000 ;
      RECT 191.620000 316.680000 234.820000 317.760000 ;
      RECT 146.620000 316.680000 189.820000 317.760000 ;
      RECT 101.620000 316.680000 144.820000 317.760000 ;
      RECT 56.620000 316.680000 99.820000 317.760000 ;
      RECT 11.620000 316.680000 54.820000 317.760000 ;
      RECT 4.860000 316.680000 9.655000 317.760000 ;
      RECT 0.000000 316.680000 2.260000 317.760000 ;
      RECT 0.000000 316.370000 548.960000 316.680000 ;
      RECT 0.000000 315.040000 550.160000 316.370000 ;
      RECT 544.900000 314.910000 550.160000 315.040000 ;
      RECT 544.900000 313.960000 548.960000 314.910000 ;
      RECT 508.620000 313.960000 542.300000 315.040000 ;
      RECT 463.620000 313.960000 506.820000 315.040000 ;
      RECT 418.620000 313.960000 461.820000 315.040000 ;
      RECT 373.620000 313.960000 416.820000 315.040000 ;
      RECT 328.620000 313.960000 371.820000 315.040000 ;
      RECT 283.620000 313.960000 326.820000 315.040000 ;
      RECT 238.620000 313.960000 281.820000 315.040000 ;
      RECT 193.620000 313.960000 236.820000 315.040000 ;
      RECT 148.620000 313.960000 191.820000 315.040000 ;
      RECT 103.620000 313.960000 146.820000 315.040000 ;
      RECT 58.620000 313.960000 101.820000 315.040000 ;
      RECT 13.620000 313.960000 56.820000 315.040000 ;
      RECT 7.860000 313.960000 11.820000 315.040000 ;
      RECT 0.000000 313.960000 5.260000 315.040000 ;
      RECT 0.000000 313.930000 548.960000 313.960000 ;
      RECT 0.000000 312.470000 550.160000 313.930000 ;
      RECT 0.000000 312.320000 548.960000 312.470000 ;
      RECT 547.900000 311.490000 548.960000 312.320000 ;
      RECT 547.900000 311.240000 550.160000 311.490000 ;
      RECT 506.620000 311.240000 545.300000 312.320000 ;
      RECT 461.620000 311.240000 504.820000 312.320000 ;
      RECT 416.620000 311.240000 459.820000 312.320000 ;
      RECT 371.620000 311.240000 414.820000 312.320000 ;
      RECT 326.620000 311.240000 369.820000 312.320000 ;
      RECT 281.620000 311.240000 324.820000 312.320000 ;
      RECT 236.620000 311.240000 279.820000 312.320000 ;
      RECT 191.620000 311.240000 234.820000 312.320000 ;
      RECT 146.620000 311.240000 189.820000 312.320000 ;
      RECT 101.620000 311.240000 144.820000 312.320000 ;
      RECT 56.620000 311.240000 99.820000 312.320000 ;
      RECT 11.620000 311.240000 54.820000 312.320000 ;
      RECT 4.860000 311.240000 9.655000 312.320000 ;
      RECT 0.000000 311.240000 2.260000 312.320000 ;
      RECT 0.000000 310.640000 550.160000 311.240000 ;
      RECT 0.000000 309.660000 548.960000 310.640000 ;
      RECT 0.000000 309.600000 550.160000 309.660000 ;
      RECT 544.900000 308.520000 550.160000 309.600000 ;
      RECT 508.620000 308.520000 542.300000 309.600000 ;
      RECT 463.620000 308.520000 506.820000 309.600000 ;
      RECT 418.620000 308.520000 461.820000 309.600000 ;
      RECT 373.620000 308.520000 416.820000 309.600000 ;
      RECT 328.620000 308.520000 371.820000 309.600000 ;
      RECT 283.620000 308.520000 326.820000 309.600000 ;
      RECT 238.620000 308.520000 281.820000 309.600000 ;
      RECT 193.620000 308.520000 236.820000 309.600000 ;
      RECT 148.620000 308.520000 191.820000 309.600000 ;
      RECT 103.620000 308.520000 146.820000 309.600000 ;
      RECT 58.620000 308.520000 101.820000 309.600000 ;
      RECT 13.620000 308.520000 56.820000 309.600000 ;
      RECT 7.860000 308.520000 11.820000 309.600000 ;
      RECT 0.000000 308.520000 5.260000 309.600000 ;
      RECT 0.000000 308.200000 550.160000 308.520000 ;
      RECT 0.000000 307.220000 548.960000 308.200000 ;
      RECT 0.000000 306.880000 550.160000 307.220000 ;
      RECT 547.900000 305.800000 550.160000 306.880000 ;
      RECT 506.620000 305.800000 545.300000 306.880000 ;
      RECT 461.620000 305.800000 504.820000 306.880000 ;
      RECT 416.620000 305.800000 459.820000 306.880000 ;
      RECT 371.620000 305.800000 414.820000 306.880000 ;
      RECT 326.620000 305.800000 369.820000 306.880000 ;
      RECT 281.620000 305.800000 324.820000 306.880000 ;
      RECT 236.620000 305.800000 279.820000 306.880000 ;
      RECT 191.620000 305.800000 234.820000 306.880000 ;
      RECT 146.620000 305.800000 189.820000 306.880000 ;
      RECT 101.620000 305.800000 144.820000 306.880000 ;
      RECT 56.620000 305.800000 99.820000 306.880000 ;
      RECT 11.620000 305.800000 54.820000 306.880000 ;
      RECT 4.860000 305.800000 9.655000 306.880000 ;
      RECT 0.000000 305.800000 2.260000 306.880000 ;
      RECT 0.000000 305.760000 550.160000 305.800000 ;
      RECT 0.000000 304.780000 548.960000 305.760000 ;
      RECT 0.000000 304.160000 550.160000 304.780000 ;
      RECT 544.900000 303.320000 550.160000 304.160000 ;
      RECT 544.900000 303.080000 548.960000 303.320000 ;
      RECT 508.620000 303.080000 542.300000 304.160000 ;
      RECT 463.620000 303.080000 506.820000 304.160000 ;
      RECT 418.620000 303.080000 461.820000 304.160000 ;
      RECT 373.620000 303.080000 416.820000 304.160000 ;
      RECT 328.620000 303.080000 371.820000 304.160000 ;
      RECT 283.620000 303.080000 326.820000 304.160000 ;
      RECT 238.620000 303.080000 281.820000 304.160000 ;
      RECT 193.620000 303.080000 236.820000 304.160000 ;
      RECT 148.620000 303.080000 191.820000 304.160000 ;
      RECT 103.620000 303.080000 146.820000 304.160000 ;
      RECT 58.620000 303.080000 101.820000 304.160000 ;
      RECT 13.620000 303.080000 56.820000 304.160000 ;
      RECT 7.860000 303.080000 11.820000 304.160000 ;
      RECT 0.000000 303.080000 5.260000 304.160000 ;
      RECT 0.000000 302.340000 548.960000 303.080000 ;
      RECT 0.000000 301.490000 550.160000 302.340000 ;
      RECT 0.000000 301.440000 548.960000 301.490000 ;
      RECT 547.900000 300.510000 548.960000 301.440000 ;
      RECT 547.900000 300.360000 550.160000 300.510000 ;
      RECT 506.620000 300.360000 545.300000 301.440000 ;
      RECT 461.620000 300.360000 504.820000 301.440000 ;
      RECT 416.620000 300.360000 459.820000 301.440000 ;
      RECT 371.620000 300.360000 414.820000 301.440000 ;
      RECT 326.620000 300.360000 369.820000 301.440000 ;
      RECT 281.620000 300.360000 324.820000 301.440000 ;
      RECT 236.620000 300.360000 279.820000 301.440000 ;
      RECT 191.620000 300.360000 234.820000 301.440000 ;
      RECT 146.620000 300.360000 189.820000 301.440000 ;
      RECT 101.620000 300.360000 144.820000 301.440000 ;
      RECT 56.620000 300.360000 99.820000 301.440000 ;
      RECT 11.620000 300.360000 54.820000 301.440000 ;
      RECT 4.860000 300.360000 9.655000 301.440000 ;
      RECT 0.000000 300.360000 2.260000 301.440000 ;
      RECT 0.000000 299.050000 550.160000 300.360000 ;
      RECT 0.000000 298.720000 548.960000 299.050000 ;
      RECT 544.900000 298.070000 548.960000 298.720000 ;
      RECT 544.900000 297.640000 550.160000 298.070000 ;
      RECT 508.620000 297.640000 542.300000 298.720000 ;
      RECT 463.620000 297.640000 506.820000 298.720000 ;
      RECT 418.620000 297.640000 461.820000 298.720000 ;
      RECT 373.620000 297.640000 416.820000 298.720000 ;
      RECT 328.620000 297.640000 371.820000 298.720000 ;
      RECT 283.620000 297.640000 326.820000 298.720000 ;
      RECT 238.620000 297.640000 281.820000 298.720000 ;
      RECT 193.620000 297.640000 236.820000 298.720000 ;
      RECT 148.620000 297.640000 191.820000 298.720000 ;
      RECT 103.620000 297.640000 146.820000 298.720000 ;
      RECT 58.620000 297.640000 101.820000 298.720000 ;
      RECT 13.620000 297.640000 56.820000 298.720000 ;
      RECT 7.860000 297.640000 11.820000 298.720000 ;
      RECT 0.000000 297.640000 5.260000 298.720000 ;
      RECT 0.000000 296.610000 550.160000 297.640000 ;
      RECT 0.000000 296.000000 548.960000 296.610000 ;
      RECT 547.900000 295.630000 548.960000 296.000000 ;
      RECT 547.900000 294.920000 550.160000 295.630000 ;
      RECT 506.620000 294.920000 545.300000 296.000000 ;
      RECT 461.620000 294.920000 504.820000 296.000000 ;
      RECT 416.620000 294.920000 459.820000 296.000000 ;
      RECT 371.620000 294.920000 414.820000 296.000000 ;
      RECT 326.620000 294.920000 369.820000 296.000000 ;
      RECT 281.620000 294.920000 324.820000 296.000000 ;
      RECT 236.620000 294.920000 279.820000 296.000000 ;
      RECT 191.620000 294.920000 234.820000 296.000000 ;
      RECT 146.620000 294.920000 189.820000 296.000000 ;
      RECT 101.620000 294.920000 144.820000 296.000000 ;
      RECT 56.620000 294.920000 99.820000 296.000000 ;
      RECT 11.620000 294.920000 54.820000 296.000000 ;
      RECT 4.860000 294.920000 9.655000 296.000000 ;
      RECT 0.000000 294.920000 2.260000 296.000000 ;
      RECT 0.000000 294.170000 550.160000 294.920000 ;
      RECT 0.000000 293.280000 548.960000 294.170000 ;
      RECT 544.900000 293.190000 548.960000 293.280000 ;
      RECT 544.900000 292.340000 550.160000 293.190000 ;
      RECT 544.900000 292.200000 548.960000 292.340000 ;
      RECT 508.620000 292.200000 542.300000 293.280000 ;
      RECT 463.620000 292.200000 506.820000 293.280000 ;
      RECT 418.620000 292.200000 461.820000 293.280000 ;
      RECT 373.620000 292.200000 416.820000 293.280000 ;
      RECT 328.620000 292.200000 371.820000 293.280000 ;
      RECT 283.620000 292.200000 326.820000 293.280000 ;
      RECT 238.620000 292.200000 281.820000 293.280000 ;
      RECT 193.620000 292.200000 236.820000 293.280000 ;
      RECT 148.620000 292.200000 191.820000 293.280000 ;
      RECT 103.620000 292.200000 146.820000 293.280000 ;
      RECT 58.620000 292.200000 101.820000 293.280000 ;
      RECT 13.620000 292.200000 56.820000 293.280000 ;
      RECT 7.860000 292.200000 11.820000 293.280000 ;
      RECT 0.000000 292.200000 5.260000 293.280000 ;
      RECT 0.000000 291.360000 548.960000 292.200000 ;
      RECT 0.000000 290.560000 550.160000 291.360000 ;
      RECT 547.900000 289.900000 550.160000 290.560000 ;
      RECT 547.900000 289.480000 548.960000 289.900000 ;
      RECT 506.620000 289.480000 545.300000 290.560000 ;
      RECT 461.620000 289.480000 504.820000 290.560000 ;
      RECT 416.620000 289.480000 459.820000 290.560000 ;
      RECT 371.620000 289.480000 414.820000 290.560000 ;
      RECT 326.620000 289.480000 369.820000 290.560000 ;
      RECT 281.620000 289.480000 324.820000 290.560000 ;
      RECT 236.620000 289.480000 279.820000 290.560000 ;
      RECT 191.620000 289.480000 234.820000 290.560000 ;
      RECT 146.620000 289.480000 189.820000 290.560000 ;
      RECT 101.620000 289.480000 144.820000 290.560000 ;
      RECT 56.620000 289.480000 99.820000 290.560000 ;
      RECT 11.620000 289.480000 54.820000 290.560000 ;
      RECT 4.860000 289.480000 9.655000 290.560000 ;
      RECT 0.000000 289.480000 2.260000 290.560000 ;
      RECT 0.000000 288.920000 548.960000 289.480000 ;
      RECT 0.000000 287.840000 550.160000 288.920000 ;
      RECT 544.900000 287.460000 550.160000 287.840000 ;
      RECT 544.900000 286.760000 548.960000 287.460000 ;
      RECT 508.620000 286.760000 542.300000 287.840000 ;
      RECT 463.620000 286.760000 506.820000 287.840000 ;
      RECT 418.620000 286.760000 461.820000 287.840000 ;
      RECT 373.620000 286.760000 416.820000 287.840000 ;
      RECT 328.620000 286.760000 371.820000 287.840000 ;
      RECT 283.620000 286.760000 326.820000 287.840000 ;
      RECT 238.620000 286.760000 281.820000 287.840000 ;
      RECT 193.620000 286.760000 236.820000 287.840000 ;
      RECT 148.620000 286.760000 191.820000 287.840000 ;
      RECT 103.620000 286.760000 146.820000 287.840000 ;
      RECT 58.620000 286.760000 101.820000 287.840000 ;
      RECT 13.620000 286.760000 56.820000 287.840000 ;
      RECT 7.860000 286.760000 11.820000 287.840000 ;
      RECT 0.000000 286.760000 5.260000 287.840000 ;
      RECT 0.000000 286.480000 548.960000 286.760000 ;
      RECT 0.000000 285.120000 550.160000 286.480000 ;
      RECT 547.900000 285.020000 550.160000 285.120000 ;
      RECT 547.900000 284.040000 548.960000 285.020000 ;
      RECT 506.620000 284.040000 545.300000 285.120000 ;
      RECT 461.620000 284.040000 504.820000 285.120000 ;
      RECT 416.620000 284.040000 459.820000 285.120000 ;
      RECT 371.620000 284.040000 414.820000 285.120000 ;
      RECT 326.620000 284.040000 369.820000 285.120000 ;
      RECT 281.620000 284.040000 324.820000 285.120000 ;
      RECT 236.620000 284.040000 279.820000 285.120000 ;
      RECT 191.620000 284.040000 234.820000 285.120000 ;
      RECT 146.620000 284.040000 189.820000 285.120000 ;
      RECT 101.620000 284.040000 144.820000 285.120000 ;
      RECT 56.620000 284.040000 99.820000 285.120000 ;
      RECT 11.620000 284.040000 54.820000 285.120000 ;
      RECT 4.860000 284.040000 9.655000 285.120000 ;
      RECT 0.000000 284.040000 2.260000 285.120000 ;
      RECT 0.000000 283.190000 550.160000 284.040000 ;
      RECT 0.000000 282.400000 548.960000 283.190000 ;
      RECT 544.900000 282.210000 548.960000 282.400000 ;
      RECT 544.900000 281.320000 550.160000 282.210000 ;
      RECT 508.620000 281.320000 542.300000 282.400000 ;
      RECT 463.620000 281.320000 506.820000 282.400000 ;
      RECT 418.620000 281.320000 461.820000 282.400000 ;
      RECT 373.620000 281.320000 416.820000 282.400000 ;
      RECT 328.620000 281.320000 371.820000 282.400000 ;
      RECT 283.620000 281.320000 326.820000 282.400000 ;
      RECT 238.620000 281.320000 281.820000 282.400000 ;
      RECT 193.620000 281.320000 236.820000 282.400000 ;
      RECT 148.620000 281.320000 191.820000 282.400000 ;
      RECT 103.620000 281.320000 146.820000 282.400000 ;
      RECT 58.620000 281.320000 101.820000 282.400000 ;
      RECT 13.620000 281.320000 56.820000 282.400000 ;
      RECT 7.860000 281.320000 11.820000 282.400000 ;
      RECT 0.000000 281.320000 5.260000 282.400000 ;
      RECT 0.000000 280.750000 550.160000 281.320000 ;
      RECT 0.000000 279.770000 548.960000 280.750000 ;
      RECT 0.000000 279.680000 550.160000 279.770000 ;
      RECT 547.900000 278.600000 550.160000 279.680000 ;
      RECT 506.620000 278.600000 545.300000 279.680000 ;
      RECT 461.620000 278.600000 504.820000 279.680000 ;
      RECT 416.620000 278.600000 459.820000 279.680000 ;
      RECT 371.620000 278.600000 414.820000 279.680000 ;
      RECT 326.620000 278.600000 369.820000 279.680000 ;
      RECT 281.620000 278.600000 324.820000 279.680000 ;
      RECT 236.620000 278.600000 279.820000 279.680000 ;
      RECT 191.620000 278.600000 234.820000 279.680000 ;
      RECT 146.620000 278.600000 189.820000 279.680000 ;
      RECT 101.620000 278.600000 144.820000 279.680000 ;
      RECT 56.620000 278.600000 99.820000 279.680000 ;
      RECT 11.620000 278.600000 54.820000 279.680000 ;
      RECT 4.860000 278.600000 9.655000 279.680000 ;
      RECT 0.000000 278.600000 2.260000 279.680000 ;
      RECT 0.000000 278.310000 550.160000 278.600000 ;
      RECT 0.000000 277.330000 548.960000 278.310000 ;
      RECT 0.000000 276.960000 550.160000 277.330000 ;
      RECT 544.900000 275.880000 550.160000 276.960000 ;
      RECT 508.620000 275.880000 542.300000 276.960000 ;
      RECT 463.620000 275.880000 506.820000 276.960000 ;
      RECT 418.620000 275.880000 461.820000 276.960000 ;
      RECT 373.620000 275.880000 416.820000 276.960000 ;
      RECT 328.620000 275.880000 371.820000 276.960000 ;
      RECT 283.620000 275.880000 326.820000 276.960000 ;
      RECT 238.620000 275.880000 281.820000 276.960000 ;
      RECT 193.620000 275.880000 236.820000 276.960000 ;
      RECT 148.620000 275.880000 191.820000 276.960000 ;
      RECT 103.620000 275.880000 146.820000 276.960000 ;
      RECT 58.620000 275.880000 101.820000 276.960000 ;
      RECT 13.620000 275.880000 56.820000 276.960000 ;
      RECT 7.860000 275.880000 11.820000 276.960000 ;
      RECT 0.000000 275.880000 5.260000 276.960000 ;
      RECT 0.000000 275.870000 550.160000 275.880000 ;
      RECT 0.000000 274.890000 548.960000 275.870000 ;
      RECT 0.000000 274.240000 550.160000 274.890000 ;
      RECT 547.900000 274.040000 550.160000 274.240000 ;
      RECT 547.900000 273.160000 548.960000 274.040000 ;
      RECT 506.620000 273.160000 545.300000 274.240000 ;
      RECT 461.620000 273.160000 504.820000 274.240000 ;
      RECT 416.620000 273.160000 459.820000 274.240000 ;
      RECT 371.620000 273.160000 414.820000 274.240000 ;
      RECT 326.620000 273.160000 369.820000 274.240000 ;
      RECT 281.620000 273.160000 324.820000 274.240000 ;
      RECT 236.620000 273.160000 279.820000 274.240000 ;
      RECT 191.620000 273.160000 234.820000 274.240000 ;
      RECT 146.620000 273.160000 189.820000 274.240000 ;
      RECT 101.620000 273.160000 144.820000 274.240000 ;
      RECT 56.620000 273.160000 99.820000 274.240000 ;
      RECT 11.620000 273.160000 54.820000 274.240000 ;
      RECT 4.860000 273.160000 9.655000 274.240000 ;
      RECT 0.000000 273.160000 2.260000 274.240000 ;
      RECT 0.000000 273.060000 548.960000 273.160000 ;
      RECT 0.000000 271.600000 550.160000 273.060000 ;
      RECT 0.000000 271.520000 548.960000 271.600000 ;
      RECT 544.900000 270.620000 548.960000 271.520000 ;
      RECT 544.900000 270.440000 550.160000 270.620000 ;
      RECT 508.620000 270.440000 542.300000 271.520000 ;
      RECT 463.620000 270.440000 506.820000 271.520000 ;
      RECT 418.620000 270.440000 461.820000 271.520000 ;
      RECT 373.620000 270.440000 416.820000 271.520000 ;
      RECT 328.620000 270.440000 371.820000 271.520000 ;
      RECT 283.620000 270.440000 326.820000 271.520000 ;
      RECT 238.620000 270.440000 281.820000 271.520000 ;
      RECT 193.620000 270.440000 236.820000 271.520000 ;
      RECT 148.620000 270.440000 191.820000 271.520000 ;
      RECT 103.620000 270.440000 146.820000 271.520000 ;
      RECT 58.620000 270.440000 101.820000 271.520000 ;
      RECT 13.620000 270.440000 56.820000 271.520000 ;
      RECT 7.860000 270.440000 11.820000 271.520000 ;
      RECT 0.000000 270.440000 5.260000 271.520000 ;
      RECT 0.000000 269.160000 550.160000 270.440000 ;
      RECT 0.000000 268.800000 548.960000 269.160000 ;
      RECT 547.900000 268.180000 548.960000 268.800000 ;
      RECT 547.900000 267.720000 550.160000 268.180000 ;
      RECT 506.620000 267.720000 545.300000 268.800000 ;
      RECT 461.620000 267.720000 504.820000 268.800000 ;
      RECT 416.620000 267.720000 459.820000 268.800000 ;
      RECT 371.620000 267.720000 414.820000 268.800000 ;
      RECT 326.620000 267.720000 369.820000 268.800000 ;
      RECT 281.620000 267.720000 324.820000 268.800000 ;
      RECT 236.620000 267.720000 279.820000 268.800000 ;
      RECT 191.620000 267.720000 234.820000 268.800000 ;
      RECT 146.620000 267.720000 189.820000 268.800000 ;
      RECT 101.620000 267.720000 144.820000 268.800000 ;
      RECT 56.620000 267.720000 99.820000 268.800000 ;
      RECT 11.620000 267.720000 54.820000 268.800000 ;
      RECT 4.860000 267.720000 9.655000 268.800000 ;
      RECT 0.000000 267.720000 2.260000 268.800000 ;
      RECT 0.000000 266.720000 550.160000 267.720000 ;
      RECT 0.000000 266.080000 548.960000 266.720000 ;
      RECT 544.900000 265.740000 548.960000 266.080000 ;
      RECT 544.900000 265.000000 550.160000 265.740000 ;
      RECT 508.620000 265.000000 542.300000 266.080000 ;
      RECT 463.620000 265.000000 506.820000 266.080000 ;
      RECT 418.620000 265.000000 461.820000 266.080000 ;
      RECT 373.620000 265.000000 416.820000 266.080000 ;
      RECT 328.620000 265.000000 371.820000 266.080000 ;
      RECT 283.620000 265.000000 326.820000 266.080000 ;
      RECT 238.620000 265.000000 281.820000 266.080000 ;
      RECT 193.620000 265.000000 236.820000 266.080000 ;
      RECT 148.620000 265.000000 191.820000 266.080000 ;
      RECT 103.620000 265.000000 146.820000 266.080000 ;
      RECT 58.620000 265.000000 101.820000 266.080000 ;
      RECT 13.620000 265.000000 56.820000 266.080000 ;
      RECT 7.860000 265.000000 11.820000 266.080000 ;
      RECT 0.000000 265.000000 5.260000 266.080000 ;
      RECT 0.000000 264.890000 550.160000 265.000000 ;
      RECT 0.000000 263.910000 548.960000 264.890000 ;
      RECT 0.000000 263.360000 550.160000 263.910000 ;
      RECT 547.900000 262.450000 550.160000 263.360000 ;
      RECT 547.900000 262.280000 548.960000 262.450000 ;
      RECT 506.620000 262.280000 545.300000 263.360000 ;
      RECT 461.620000 262.280000 504.820000 263.360000 ;
      RECT 416.620000 262.280000 459.820000 263.360000 ;
      RECT 371.620000 262.280000 414.820000 263.360000 ;
      RECT 326.620000 262.280000 369.820000 263.360000 ;
      RECT 281.620000 262.280000 324.820000 263.360000 ;
      RECT 236.620000 262.280000 279.820000 263.360000 ;
      RECT 191.620000 262.280000 234.820000 263.360000 ;
      RECT 146.620000 262.280000 189.820000 263.360000 ;
      RECT 101.620000 262.280000 144.820000 263.360000 ;
      RECT 56.620000 262.280000 99.820000 263.360000 ;
      RECT 11.620000 262.280000 54.820000 263.360000 ;
      RECT 4.860000 262.280000 9.655000 263.360000 ;
      RECT 0.000000 262.280000 2.260000 263.360000 ;
      RECT 0.000000 261.470000 548.960000 262.280000 ;
      RECT 0.000000 260.640000 550.160000 261.470000 ;
      RECT 544.900000 260.010000 550.160000 260.640000 ;
      RECT 544.900000 259.560000 548.960000 260.010000 ;
      RECT 508.620000 259.560000 542.300000 260.640000 ;
      RECT 463.620000 259.560000 506.820000 260.640000 ;
      RECT 418.620000 259.560000 461.820000 260.640000 ;
      RECT 373.620000 259.560000 416.820000 260.640000 ;
      RECT 328.620000 259.560000 371.820000 260.640000 ;
      RECT 283.620000 259.560000 326.820000 260.640000 ;
      RECT 238.620000 259.560000 281.820000 260.640000 ;
      RECT 193.620000 259.560000 236.820000 260.640000 ;
      RECT 148.620000 259.560000 191.820000 260.640000 ;
      RECT 103.620000 259.560000 146.820000 260.640000 ;
      RECT 58.620000 259.560000 101.820000 260.640000 ;
      RECT 13.620000 259.560000 56.820000 260.640000 ;
      RECT 7.860000 259.560000 11.820000 260.640000 ;
      RECT 0.000000 259.560000 5.260000 260.640000 ;
      RECT 0.000000 259.030000 548.960000 259.560000 ;
      RECT 0.000000 257.920000 550.160000 259.030000 ;
      RECT 547.900000 257.570000 550.160000 257.920000 ;
      RECT 547.900000 256.840000 548.960000 257.570000 ;
      RECT 506.620000 256.840000 545.300000 257.920000 ;
      RECT 461.620000 256.840000 504.820000 257.920000 ;
      RECT 416.620000 256.840000 459.820000 257.920000 ;
      RECT 371.620000 256.840000 414.820000 257.920000 ;
      RECT 326.620000 256.840000 369.820000 257.920000 ;
      RECT 281.620000 256.840000 324.820000 257.920000 ;
      RECT 236.620000 256.840000 279.820000 257.920000 ;
      RECT 191.620000 256.840000 234.820000 257.920000 ;
      RECT 146.620000 256.840000 189.820000 257.920000 ;
      RECT 101.620000 256.840000 144.820000 257.920000 ;
      RECT 56.620000 256.840000 99.820000 257.920000 ;
      RECT 11.620000 256.840000 54.820000 257.920000 ;
      RECT 4.860000 256.840000 9.655000 257.920000 ;
      RECT 0.000000 256.840000 2.260000 257.920000 ;
      RECT 0.000000 256.590000 548.960000 256.840000 ;
      RECT 0.000000 255.740000 550.160000 256.590000 ;
      RECT 0.000000 255.200000 548.960000 255.740000 ;
      RECT 544.900000 254.760000 548.960000 255.200000 ;
      RECT 544.900000 254.120000 550.160000 254.760000 ;
      RECT 508.620000 254.120000 542.300000 255.200000 ;
      RECT 463.620000 254.120000 506.820000 255.200000 ;
      RECT 418.620000 254.120000 461.820000 255.200000 ;
      RECT 373.620000 254.120000 416.820000 255.200000 ;
      RECT 328.620000 254.120000 371.820000 255.200000 ;
      RECT 283.620000 254.120000 326.820000 255.200000 ;
      RECT 238.620000 254.120000 281.820000 255.200000 ;
      RECT 193.620000 254.120000 236.820000 255.200000 ;
      RECT 148.620000 254.120000 191.820000 255.200000 ;
      RECT 103.620000 254.120000 146.820000 255.200000 ;
      RECT 58.620000 254.120000 101.820000 255.200000 ;
      RECT 13.620000 254.120000 56.820000 255.200000 ;
      RECT 7.860000 254.120000 11.820000 255.200000 ;
      RECT 0.000000 254.120000 5.260000 255.200000 ;
      RECT 0.000000 253.300000 550.160000 254.120000 ;
      RECT 0.000000 252.480000 548.960000 253.300000 ;
      RECT 547.900000 252.320000 548.960000 252.480000 ;
      RECT 547.900000 251.400000 550.160000 252.320000 ;
      RECT 506.620000 251.400000 545.300000 252.480000 ;
      RECT 461.620000 251.400000 504.820000 252.480000 ;
      RECT 416.620000 251.400000 459.820000 252.480000 ;
      RECT 371.620000 251.400000 414.820000 252.480000 ;
      RECT 326.620000 251.400000 369.820000 252.480000 ;
      RECT 281.620000 251.400000 324.820000 252.480000 ;
      RECT 236.620000 251.400000 279.820000 252.480000 ;
      RECT 191.620000 251.400000 234.820000 252.480000 ;
      RECT 146.620000 251.400000 189.820000 252.480000 ;
      RECT 101.620000 251.400000 144.820000 252.480000 ;
      RECT 56.620000 251.400000 99.820000 252.480000 ;
      RECT 11.620000 251.400000 54.820000 252.480000 ;
      RECT 4.860000 251.400000 9.655000 252.480000 ;
      RECT 0.000000 251.400000 2.260000 252.480000 ;
      RECT 0.000000 250.860000 550.160000 251.400000 ;
      RECT 0.000000 249.880000 548.960000 250.860000 ;
      RECT 0.000000 249.760000 550.160000 249.880000 ;
      RECT 544.900000 248.680000 550.160000 249.760000 ;
      RECT 508.620000 248.680000 542.300000 249.760000 ;
      RECT 463.620000 248.680000 506.820000 249.760000 ;
      RECT 418.620000 248.680000 461.820000 249.760000 ;
      RECT 373.620000 248.680000 416.820000 249.760000 ;
      RECT 328.620000 248.680000 371.820000 249.760000 ;
      RECT 283.620000 248.680000 326.820000 249.760000 ;
      RECT 238.620000 248.680000 281.820000 249.760000 ;
      RECT 193.620000 248.680000 236.820000 249.760000 ;
      RECT 148.620000 248.680000 191.820000 249.760000 ;
      RECT 103.620000 248.680000 146.820000 249.760000 ;
      RECT 58.620000 248.680000 101.820000 249.760000 ;
      RECT 13.620000 248.680000 56.820000 249.760000 ;
      RECT 7.860000 248.680000 11.820000 249.760000 ;
      RECT 0.000000 248.680000 5.260000 249.760000 ;
      RECT 0.000000 248.420000 550.160000 248.680000 ;
      RECT 0.000000 247.440000 548.960000 248.420000 ;
      RECT 0.000000 247.040000 550.160000 247.440000 ;
      RECT 547.900000 246.590000 550.160000 247.040000 ;
      RECT 547.900000 245.960000 548.960000 246.590000 ;
      RECT 506.620000 245.960000 545.300000 247.040000 ;
      RECT 461.620000 245.960000 504.820000 247.040000 ;
      RECT 416.620000 245.960000 459.820000 247.040000 ;
      RECT 371.620000 245.960000 414.820000 247.040000 ;
      RECT 326.620000 245.960000 369.820000 247.040000 ;
      RECT 281.620000 245.960000 324.820000 247.040000 ;
      RECT 236.620000 245.960000 279.820000 247.040000 ;
      RECT 191.620000 245.960000 234.820000 247.040000 ;
      RECT 146.620000 245.960000 189.820000 247.040000 ;
      RECT 101.620000 245.960000 144.820000 247.040000 ;
      RECT 56.620000 245.960000 99.820000 247.040000 ;
      RECT 11.620000 245.960000 54.820000 247.040000 ;
      RECT 4.860000 245.960000 9.655000 247.040000 ;
      RECT 0.000000 245.960000 2.260000 247.040000 ;
      RECT 0.000000 245.610000 548.960000 245.960000 ;
      RECT 0.000000 244.320000 550.160000 245.610000 ;
      RECT 544.900000 244.150000 550.160000 244.320000 ;
      RECT 544.900000 243.240000 548.960000 244.150000 ;
      RECT 508.620000 243.240000 542.300000 244.320000 ;
      RECT 463.620000 243.240000 506.820000 244.320000 ;
      RECT 418.620000 243.240000 461.820000 244.320000 ;
      RECT 373.620000 243.240000 416.820000 244.320000 ;
      RECT 328.620000 243.240000 371.820000 244.320000 ;
      RECT 283.620000 243.240000 326.820000 244.320000 ;
      RECT 238.620000 243.240000 281.820000 244.320000 ;
      RECT 193.620000 243.240000 236.820000 244.320000 ;
      RECT 148.620000 243.240000 191.820000 244.320000 ;
      RECT 103.620000 243.240000 146.820000 244.320000 ;
      RECT 58.620000 243.240000 101.820000 244.320000 ;
      RECT 13.620000 243.240000 56.820000 244.320000 ;
      RECT 7.860000 243.240000 11.820000 244.320000 ;
      RECT 0.000000 243.240000 5.260000 244.320000 ;
      RECT 0.000000 243.170000 548.960000 243.240000 ;
      RECT 0.000000 241.710000 550.160000 243.170000 ;
      RECT 0.000000 241.600000 548.960000 241.710000 ;
      RECT 547.900000 240.730000 548.960000 241.600000 ;
      RECT 547.900000 240.520000 550.160000 240.730000 ;
      RECT 506.620000 240.520000 545.300000 241.600000 ;
      RECT 461.620000 240.520000 504.820000 241.600000 ;
      RECT 416.620000 240.520000 459.820000 241.600000 ;
      RECT 371.620000 240.520000 414.820000 241.600000 ;
      RECT 326.620000 240.520000 369.820000 241.600000 ;
      RECT 281.620000 240.520000 324.820000 241.600000 ;
      RECT 236.620000 240.520000 279.820000 241.600000 ;
      RECT 191.620000 240.520000 234.820000 241.600000 ;
      RECT 146.620000 240.520000 189.820000 241.600000 ;
      RECT 101.620000 240.520000 144.820000 241.600000 ;
      RECT 56.620000 240.520000 99.820000 241.600000 ;
      RECT 11.620000 240.520000 54.820000 241.600000 ;
      RECT 4.860000 240.520000 9.655000 241.600000 ;
      RECT 0.000000 240.520000 2.260000 241.600000 ;
      RECT 0.000000 239.270000 550.160000 240.520000 ;
      RECT 0.000000 238.880000 548.960000 239.270000 ;
      RECT 544.900000 238.290000 548.960000 238.880000 ;
      RECT 544.900000 237.800000 550.160000 238.290000 ;
      RECT 508.620000 237.800000 542.300000 238.880000 ;
      RECT 463.620000 237.800000 506.820000 238.880000 ;
      RECT 418.620000 237.800000 461.820000 238.880000 ;
      RECT 373.620000 237.800000 416.820000 238.880000 ;
      RECT 328.620000 237.800000 371.820000 238.880000 ;
      RECT 283.620000 237.800000 326.820000 238.880000 ;
      RECT 238.620000 237.800000 281.820000 238.880000 ;
      RECT 193.620000 237.800000 236.820000 238.880000 ;
      RECT 148.620000 237.800000 191.820000 238.880000 ;
      RECT 103.620000 237.800000 146.820000 238.880000 ;
      RECT 58.620000 237.800000 101.820000 238.880000 ;
      RECT 13.620000 237.800000 56.820000 238.880000 ;
      RECT 7.860000 237.800000 11.820000 238.880000 ;
      RECT 0.000000 237.800000 5.260000 238.880000 ;
      RECT 0.000000 236.830000 550.160000 237.800000 ;
      RECT 0.000000 236.160000 548.960000 236.830000 ;
      RECT 547.900000 235.850000 548.960000 236.160000 ;
      RECT 547.900000 235.080000 550.160000 235.850000 ;
      RECT 506.620000 235.080000 545.300000 236.160000 ;
      RECT 461.620000 235.080000 504.820000 236.160000 ;
      RECT 416.620000 235.080000 459.820000 236.160000 ;
      RECT 371.620000 235.080000 414.820000 236.160000 ;
      RECT 326.620000 235.080000 369.820000 236.160000 ;
      RECT 281.620000 235.080000 324.820000 236.160000 ;
      RECT 236.620000 235.080000 279.820000 236.160000 ;
      RECT 191.620000 235.080000 234.820000 236.160000 ;
      RECT 146.620000 235.080000 189.820000 236.160000 ;
      RECT 101.620000 235.080000 144.820000 236.160000 ;
      RECT 56.620000 235.080000 99.820000 236.160000 ;
      RECT 11.620000 235.080000 54.820000 236.160000 ;
      RECT 4.860000 235.080000 9.655000 236.160000 ;
      RECT 0.000000 235.080000 2.260000 236.160000 ;
      RECT 0.000000 235.000000 550.160000 235.080000 ;
      RECT 0.000000 234.020000 548.960000 235.000000 ;
      RECT 0.000000 233.440000 550.160000 234.020000 ;
      RECT 544.900000 232.560000 550.160000 233.440000 ;
      RECT 544.900000 232.360000 548.960000 232.560000 ;
      RECT 508.620000 232.360000 542.300000 233.440000 ;
      RECT 463.620000 232.360000 506.820000 233.440000 ;
      RECT 418.620000 232.360000 461.820000 233.440000 ;
      RECT 373.620000 232.360000 416.820000 233.440000 ;
      RECT 328.620000 232.360000 371.820000 233.440000 ;
      RECT 283.620000 232.360000 326.820000 233.440000 ;
      RECT 238.620000 232.360000 281.820000 233.440000 ;
      RECT 193.620000 232.360000 236.820000 233.440000 ;
      RECT 148.620000 232.360000 191.820000 233.440000 ;
      RECT 103.620000 232.360000 146.820000 233.440000 ;
      RECT 58.620000 232.360000 101.820000 233.440000 ;
      RECT 13.620000 232.360000 56.820000 233.440000 ;
      RECT 7.860000 232.360000 11.820000 233.440000 ;
      RECT 0.000000 232.360000 5.260000 233.440000 ;
      RECT 0.000000 231.580000 548.960000 232.360000 ;
      RECT 0.000000 230.720000 550.160000 231.580000 ;
      RECT 547.900000 230.120000 550.160000 230.720000 ;
      RECT 547.900000 229.640000 548.960000 230.120000 ;
      RECT 506.620000 229.640000 545.300000 230.720000 ;
      RECT 461.620000 229.640000 504.820000 230.720000 ;
      RECT 416.620000 229.640000 459.820000 230.720000 ;
      RECT 371.620000 229.640000 414.820000 230.720000 ;
      RECT 326.620000 229.640000 369.820000 230.720000 ;
      RECT 281.620000 229.640000 324.820000 230.720000 ;
      RECT 236.620000 229.640000 279.820000 230.720000 ;
      RECT 191.620000 229.640000 234.820000 230.720000 ;
      RECT 146.620000 229.640000 189.820000 230.720000 ;
      RECT 101.620000 229.640000 144.820000 230.720000 ;
      RECT 56.620000 229.640000 99.820000 230.720000 ;
      RECT 11.620000 229.640000 54.820000 230.720000 ;
      RECT 4.860000 229.640000 9.655000 230.720000 ;
      RECT 0.000000 229.640000 2.260000 230.720000 ;
      RECT 0.000000 229.140000 548.960000 229.640000 ;
      RECT 0.000000 228.000000 550.160000 229.140000 ;
      RECT 544.900000 227.680000 550.160000 228.000000 ;
      RECT 544.900000 226.920000 548.960000 227.680000 ;
      RECT 508.620000 226.920000 542.300000 228.000000 ;
      RECT 463.620000 226.920000 506.820000 228.000000 ;
      RECT 418.620000 226.920000 461.820000 228.000000 ;
      RECT 373.620000 226.920000 416.820000 228.000000 ;
      RECT 328.620000 226.920000 371.820000 228.000000 ;
      RECT 283.620000 226.920000 326.820000 228.000000 ;
      RECT 238.620000 226.920000 281.820000 228.000000 ;
      RECT 193.620000 226.920000 236.820000 228.000000 ;
      RECT 148.620000 226.920000 191.820000 228.000000 ;
      RECT 103.620000 226.920000 146.820000 228.000000 ;
      RECT 58.620000 226.920000 101.820000 228.000000 ;
      RECT 13.620000 226.920000 56.820000 228.000000 ;
      RECT 7.860000 226.920000 11.820000 228.000000 ;
      RECT 0.000000 226.920000 5.260000 228.000000 ;
      RECT 0.000000 226.700000 548.960000 226.920000 ;
      RECT 0.000000 225.850000 550.160000 226.700000 ;
      RECT 0.000000 225.280000 548.960000 225.850000 ;
      RECT 547.900000 224.870000 548.960000 225.280000 ;
      RECT 547.900000 224.200000 550.160000 224.870000 ;
      RECT 506.620000 224.200000 545.300000 225.280000 ;
      RECT 461.620000 224.200000 504.820000 225.280000 ;
      RECT 416.620000 224.200000 459.820000 225.280000 ;
      RECT 371.620000 224.200000 414.820000 225.280000 ;
      RECT 326.620000 224.200000 369.820000 225.280000 ;
      RECT 281.620000 224.200000 324.820000 225.280000 ;
      RECT 236.620000 224.200000 279.820000 225.280000 ;
      RECT 191.620000 224.200000 234.820000 225.280000 ;
      RECT 146.620000 224.200000 189.820000 225.280000 ;
      RECT 101.620000 224.200000 144.820000 225.280000 ;
      RECT 56.620000 224.200000 99.820000 225.280000 ;
      RECT 11.620000 224.200000 54.820000 225.280000 ;
      RECT 4.860000 224.200000 9.655000 225.280000 ;
      RECT 0.000000 224.200000 2.260000 225.280000 ;
      RECT 0.000000 223.410000 550.160000 224.200000 ;
      RECT 0.000000 222.560000 548.960000 223.410000 ;
      RECT 544.900000 222.430000 548.960000 222.560000 ;
      RECT 544.900000 221.480000 550.160000 222.430000 ;
      RECT 508.620000 221.480000 542.300000 222.560000 ;
      RECT 463.620000 221.480000 506.820000 222.560000 ;
      RECT 418.620000 221.480000 461.820000 222.560000 ;
      RECT 373.620000 221.480000 416.820000 222.560000 ;
      RECT 328.620000 221.480000 371.820000 222.560000 ;
      RECT 283.620000 221.480000 326.820000 222.560000 ;
      RECT 238.620000 221.480000 281.820000 222.560000 ;
      RECT 193.620000 221.480000 236.820000 222.560000 ;
      RECT 148.620000 221.480000 191.820000 222.560000 ;
      RECT 103.620000 221.480000 146.820000 222.560000 ;
      RECT 58.620000 221.480000 101.820000 222.560000 ;
      RECT 13.620000 221.480000 56.820000 222.560000 ;
      RECT 7.860000 221.480000 11.820000 222.560000 ;
      RECT 0.000000 221.480000 5.260000 222.560000 ;
      RECT 0.000000 220.970000 550.160000 221.480000 ;
      RECT 0.000000 219.990000 548.960000 220.970000 ;
      RECT 0.000000 219.840000 550.160000 219.990000 ;
      RECT 547.900000 218.760000 550.160000 219.840000 ;
      RECT 506.620000 218.760000 545.300000 219.840000 ;
      RECT 461.620000 218.760000 504.820000 219.840000 ;
      RECT 416.620000 218.760000 459.820000 219.840000 ;
      RECT 371.620000 218.760000 414.820000 219.840000 ;
      RECT 326.620000 218.760000 369.820000 219.840000 ;
      RECT 281.620000 218.760000 324.820000 219.840000 ;
      RECT 236.620000 218.760000 279.820000 219.840000 ;
      RECT 191.620000 218.760000 234.820000 219.840000 ;
      RECT 146.620000 218.760000 189.820000 219.840000 ;
      RECT 101.620000 218.760000 144.820000 219.840000 ;
      RECT 56.620000 218.760000 99.820000 219.840000 ;
      RECT 11.620000 218.760000 54.820000 219.840000 ;
      RECT 4.860000 218.760000 9.655000 219.840000 ;
      RECT 0.000000 218.760000 2.260000 219.840000 ;
      RECT 0.000000 218.530000 550.160000 218.760000 ;
      RECT 0.000000 217.550000 548.960000 218.530000 ;
      RECT 0.000000 217.120000 550.160000 217.550000 ;
      RECT 544.900000 216.700000 550.160000 217.120000 ;
      RECT 544.900000 216.040000 548.960000 216.700000 ;
      RECT 508.620000 216.040000 542.300000 217.120000 ;
      RECT 463.620000 216.040000 506.820000 217.120000 ;
      RECT 418.620000 216.040000 461.820000 217.120000 ;
      RECT 373.620000 216.040000 416.820000 217.120000 ;
      RECT 328.620000 216.040000 371.820000 217.120000 ;
      RECT 283.620000 216.040000 326.820000 217.120000 ;
      RECT 238.620000 216.040000 281.820000 217.120000 ;
      RECT 193.620000 216.040000 236.820000 217.120000 ;
      RECT 148.620000 216.040000 191.820000 217.120000 ;
      RECT 103.620000 216.040000 146.820000 217.120000 ;
      RECT 58.620000 216.040000 101.820000 217.120000 ;
      RECT 13.620000 216.040000 56.820000 217.120000 ;
      RECT 7.860000 216.040000 11.820000 217.120000 ;
      RECT 0.000000 216.040000 5.260000 217.120000 ;
      RECT 0.000000 215.720000 548.960000 216.040000 ;
      RECT 0.000000 214.400000 550.160000 215.720000 ;
      RECT 547.900000 214.260000 550.160000 214.400000 ;
      RECT 547.900000 213.320000 548.960000 214.260000 ;
      RECT 506.620000 213.320000 545.300000 214.400000 ;
      RECT 461.620000 213.320000 504.820000 214.400000 ;
      RECT 416.620000 213.320000 459.820000 214.400000 ;
      RECT 371.620000 213.320000 414.820000 214.400000 ;
      RECT 326.620000 213.320000 369.820000 214.400000 ;
      RECT 281.620000 213.320000 324.820000 214.400000 ;
      RECT 236.620000 213.320000 279.820000 214.400000 ;
      RECT 191.620000 213.320000 234.820000 214.400000 ;
      RECT 146.620000 213.320000 189.820000 214.400000 ;
      RECT 101.620000 213.320000 144.820000 214.400000 ;
      RECT 56.620000 213.320000 99.820000 214.400000 ;
      RECT 11.620000 213.320000 54.820000 214.400000 ;
      RECT 4.860000 213.320000 9.655000 214.400000 ;
      RECT 0.000000 213.320000 2.260000 214.400000 ;
      RECT 0.000000 213.280000 548.960000 213.320000 ;
      RECT 0.000000 211.820000 550.160000 213.280000 ;
      RECT 0.000000 211.680000 548.960000 211.820000 ;
      RECT 544.900000 210.840000 548.960000 211.680000 ;
      RECT 544.900000 210.600000 550.160000 210.840000 ;
      RECT 508.620000 210.600000 542.300000 211.680000 ;
      RECT 463.620000 210.600000 506.820000 211.680000 ;
      RECT 418.620000 210.600000 461.820000 211.680000 ;
      RECT 373.620000 210.600000 416.820000 211.680000 ;
      RECT 328.620000 210.600000 371.820000 211.680000 ;
      RECT 283.620000 210.600000 326.820000 211.680000 ;
      RECT 238.620000 210.600000 281.820000 211.680000 ;
      RECT 193.620000 210.600000 236.820000 211.680000 ;
      RECT 148.620000 210.600000 191.820000 211.680000 ;
      RECT 103.620000 210.600000 146.820000 211.680000 ;
      RECT 58.620000 210.600000 101.820000 211.680000 ;
      RECT 13.620000 210.600000 56.820000 211.680000 ;
      RECT 7.860000 210.600000 11.820000 211.680000 ;
      RECT 0.000000 210.600000 5.260000 211.680000 ;
      RECT 0.000000 209.380000 550.160000 210.600000 ;
      RECT 0.000000 208.960000 548.960000 209.380000 ;
      RECT 547.900000 208.400000 548.960000 208.960000 ;
      RECT 547.900000 207.880000 550.160000 208.400000 ;
      RECT 506.620000 207.880000 545.300000 208.960000 ;
      RECT 461.620000 207.880000 504.820000 208.960000 ;
      RECT 416.620000 207.880000 459.820000 208.960000 ;
      RECT 371.620000 207.880000 414.820000 208.960000 ;
      RECT 326.620000 207.880000 369.820000 208.960000 ;
      RECT 281.620000 207.880000 324.820000 208.960000 ;
      RECT 236.620000 207.880000 279.820000 208.960000 ;
      RECT 191.620000 207.880000 234.820000 208.960000 ;
      RECT 146.620000 207.880000 189.820000 208.960000 ;
      RECT 101.620000 207.880000 144.820000 208.960000 ;
      RECT 56.620000 207.880000 99.820000 208.960000 ;
      RECT 11.620000 207.880000 54.820000 208.960000 ;
      RECT 4.860000 207.880000 9.655000 208.960000 ;
      RECT 0.000000 207.880000 2.260000 208.960000 ;
      RECT 0.000000 207.550000 550.160000 207.880000 ;
      RECT 0.000000 206.570000 548.960000 207.550000 ;
      RECT 0.000000 206.240000 550.160000 206.570000 ;
      RECT 544.900000 205.160000 550.160000 206.240000 ;
      RECT 508.620000 205.160000 542.300000 206.240000 ;
      RECT 463.620000 205.160000 506.820000 206.240000 ;
      RECT 418.620000 205.160000 461.820000 206.240000 ;
      RECT 373.620000 205.160000 416.820000 206.240000 ;
      RECT 328.620000 205.160000 371.820000 206.240000 ;
      RECT 283.620000 205.160000 326.820000 206.240000 ;
      RECT 238.620000 205.160000 281.820000 206.240000 ;
      RECT 193.620000 205.160000 236.820000 206.240000 ;
      RECT 148.620000 205.160000 191.820000 206.240000 ;
      RECT 103.620000 205.160000 146.820000 206.240000 ;
      RECT 58.620000 205.160000 101.820000 206.240000 ;
      RECT 13.620000 205.160000 56.820000 206.240000 ;
      RECT 7.860000 205.160000 11.820000 206.240000 ;
      RECT 0.000000 205.160000 5.260000 206.240000 ;
      RECT 0.000000 205.110000 550.160000 205.160000 ;
      RECT 0.000000 204.130000 548.960000 205.110000 ;
      RECT 0.000000 203.520000 550.160000 204.130000 ;
      RECT 547.900000 202.670000 550.160000 203.520000 ;
      RECT 547.900000 202.440000 548.960000 202.670000 ;
      RECT 506.620000 202.440000 545.300000 203.520000 ;
      RECT 461.620000 202.440000 504.820000 203.520000 ;
      RECT 416.620000 202.440000 459.820000 203.520000 ;
      RECT 371.620000 202.440000 414.820000 203.520000 ;
      RECT 326.620000 202.440000 369.820000 203.520000 ;
      RECT 281.620000 202.440000 324.820000 203.520000 ;
      RECT 236.620000 202.440000 279.820000 203.520000 ;
      RECT 191.620000 202.440000 234.820000 203.520000 ;
      RECT 146.620000 202.440000 189.820000 203.520000 ;
      RECT 101.620000 202.440000 144.820000 203.520000 ;
      RECT 56.620000 202.440000 99.820000 203.520000 ;
      RECT 11.620000 202.440000 54.820000 203.520000 ;
      RECT 4.860000 202.440000 9.655000 203.520000 ;
      RECT 0.000000 202.440000 2.260000 203.520000 ;
      RECT 0.000000 201.690000 548.960000 202.440000 ;
      RECT 0.000000 200.800000 550.160000 201.690000 ;
      RECT 544.900000 200.230000 550.160000 200.800000 ;
      RECT 544.900000 199.720000 548.960000 200.230000 ;
      RECT 508.620000 199.720000 542.300000 200.800000 ;
      RECT 463.620000 199.720000 506.820000 200.800000 ;
      RECT 418.620000 199.720000 461.820000 200.800000 ;
      RECT 373.620000 199.720000 416.820000 200.800000 ;
      RECT 328.620000 199.720000 371.820000 200.800000 ;
      RECT 283.620000 199.720000 326.820000 200.800000 ;
      RECT 238.620000 199.720000 281.820000 200.800000 ;
      RECT 193.620000 199.720000 236.820000 200.800000 ;
      RECT 148.620000 199.720000 191.820000 200.800000 ;
      RECT 103.620000 199.720000 146.820000 200.800000 ;
      RECT 58.620000 199.720000 101.820000 200.800000 ;
      RECT 13.620000 199.720000 56.820000 200.800000 ;
      RECT 7.860000 199.720000 11.820000 200.800000 ;
      RECT 0.000000 199.720000 5.260000 200.800000 ;
      RECT 0.000000 199.250000 548.960000 199.720000 ;
      RECT 0.000000 198.400000 550.160000 199.250000 ;
      RECT 0.000000 198.080000 548.960000 198.400000 ;
      RECT 547.900000 197.420000 548.960000 198.080000 ;
      RECT 547.900000 197.000000 550.160000 197.420000 ;
      RECT 506.620000 197.000000 545.300000 198.080000 ;
      RECT 461.620000 197.000000 504.820000 198.080000 ;
      RECT 416.620000 197.000000 459.820000 198.080000 ;
      RECT 371.620000 197.000000 414.820000 198.080000 ;
      RECT 326.620000 197.000000 369.820000 198.080000 ;
      RECT 281.620000 197.000000 324.820000 198.080000 ;
      RECT 236.620000 197.000000 279.820000 198.080000 ;
      RECT 191.620000 197.000000 234.820000 198.080000 ;
      RECT 146.620000 197.000000 189.820000 198.080000 ;
      RECT 101.620000 197.000000 144.820000 198.080000 ;
      RECT 56.620000 197.000000 99.820000 198.080000 ;
      RECT 11.620000 197.000000 54.820000 198.080000 ;
      RECT 4.860000 197.000000 9.655000 198.080000 ;
      RECT 0.000000 197.000000 2.260000 198.080000 ;
      RECT 0.000000 195.960000 550.160000 197.000000 ;
      RECT 0.000000 195.360000 548.960000 195.960000 ;
      RECT 544.900000 194.980000 548.960000 195.360000 ;
      RECT 544.900000 194.280000 550.160000 194.980000 ;
      RECT 508.620000 194.280000 542.300000 195.360000 ;
      RECT 463.620000 194.280000 506.820000 195.360000 ;
      RECT 418.620000 194.280000 461.820000 195.360000 ;
      RECT 373.620000 194.280000 416.820000 195.360000 ;
      RECT 328.620000 194.280000 371.820000 195.360000 ;
      RECT 283.620000 194.280000 326.820000 195.360000 ;
      RECT 238.620000 194.280000 281.820000 195.360000 ;
      RECT 193.620000 194.280000 236.820000 195.360000 ;
      RECT 148.620000 194.280000 191.820000 195.360000 ;
      RECT 103.620000 194.280000 146.820000 195.360000 ;
      RECT 58.620000 194.280000 101.820000 195.360000 ;
      RECT 13.620000 194.280000 56.820000 195.360000 ;
      RECT 7.860000 194.280000 11.820000 195.360000 ;
      RECT 0.000000 194.280000 5.260000 195.360000 ;
      RECT 0.000000 193.520000 550.160000 194.280000 ;
      RECT 0.000000 192.640000 548.960000 193.520000 ;
      RECT 547.900000 192.540000 548.960000 192.640000 ;
      RECT 547.900000 191.560000 550.160000 192.540000 ;
      RECT 506.620000 191.560000 545.300000 192.640000 ;
      RECT 461.620000 191.560000 504.820000 192.640000 ;
      RECT 416.620000 191.560000 459.820000 192.640000 ;
      RECT 371.620000 191.560000 414.820000 192.640000 ;
      RECT 326.620000 191.560000 369.820000 192.640000 ;
      RECT 281.620000 191.560000 324.820000 192.640000 ;
      RECT 236.620000 191.560000 279.820000 192.640000 ;
      RECT 191.620000 191.560000 234.820000 192.640000 ;
      RECT 146.620000 191.560000 189.820000 192.640000 ;
      RECT 101.620000 191.560000 144.820000 192.640000 ;
      RECT 56.620000 191.560000 99.820000 192.640000 ;
      RECT 11.620000 191.560000 54.820000 192.640000 ;
      RECT 4.860000 191.560000 9.655000 192.640000 ;
      RECT 0.000000 191.560000 2.260000 192.640000 ;
      RECT 0.000000 191.080000 550.160000 191.560000 ;
      RECT 0.000000 190.100000 548.960000 191.080000 ;
      RECT 0.000000 189.920000 550.160000 190.100000 ;
      RECT 544.900000 189.250000 550.160000 189.920000 ;
      RECT 544.900000 188.840000 548.960000 189.250000 ;
      RECT 508.620000 188.840000 542.300000 189.920000 ;
      RECT 463.620000 188.840000 506.820000 189.920000 ;
      RECT 418.620000 188.840000 461.820000 189.920000 ;
      RECT 373.620000 188.840000 416.820000 189.920000 ;
      RECT 328.620000 188.840000 371.820000 189.920000 ;
      RECT 283.620000 188.840000 326.820000 189.920000 ;
      RECT 238.620000 188.840000 281.820000 189.920000 ;
      RECT 193.620000 188.840000 236.820000 189.920000 ;
      RECT 148.620000 188.840000 191.820000 189.920000 ;
      RECT 103.620000 188.840000 146.820000 189.920000 ;
      RECT 58.620000 188.840000 101.820000 189.920000 ;
      RECT 13.620000 188.840000 56.820000 189.920000 ;
      RECT 7.860000 188.840000 11.820000 189.920000 ;
      RECT 0.000000 188.840000 5.260000 189.920000 ;
      RECT 0.000000 188.270000 548.960000 188.840000 ;
      RECT 0.000000 187.200000 550.160000 188.270000 ;
      RECT 547.900000 186.810000 550.160000 187.200000 ;
      RECT 547.900000 186.120000 548.960000 186.810000 ;
      RECT 506.620000 186.120000 545.300000 187.200000 ;
      RECT 461.620000 186.120000 504.820000 187.200000 ;
      RECT 416.620000 186.120000 459.820000 187.200000 ;
      RECT 371.620000 186.120000 414.820000 187.200000 ;
      RECT 326.620000 186.120000 369.820000 187.200000 ;
      RECT 281.620000 186.120000 324.820000 187.200000 ;
      RECT 236.620000 186.120000 279.820000 187.200000 ;
      RECT 191.620000 186.120000 234.820000 187.200000 ;
      RECT 146.620000 186.120000 189.820000 187.200000 ;
      RECT 101.620000 186.120000 144.820000 187.200000 ;
      RECT 56.620000 186.120000 99.820000 187.200000 ;
      RECT 11.620000 186.120000 54.820000 187.200000 ;
      RECT 4.860000 186.120000 9.655000 187.200000 ;
      RECT 0.000000 186.120000 2.260000 187.200000 ;
      RECT 0.000000 185.830000 548.960000 186.120000 ;
      RECT 0.000000 184.480000 550.160000 185.830000 ;
      RECT 544.900000 184.370000 550.160000 184.480000 ;
      RECT 544.900000 183.400000 548.960000 184.370000 ;
      RECT 508.620000 183.400000 542.300000 184.480000 ;
      RECT 463.620000 183.400000 506.820000 184.480000 ;
      RECT 418.620000 183.400000 461.820000 184.480000 ;
      RECT 373.620000 183.400000 416.820000 184.480000 ;
      RECT 328.620000 183.400000 371.820000 184.480000 ;
      RECT 283.620000 183.400000 326.820000 184.480000 ;
      RECT 238.620000 183.400000 281.820000 184.480000 ;
      RECT 193.620000 183.400000 236.820000 184.480000 ;
      RECT 148.620000 183.400000 191.820000 184.480000 ;
      RECT 103.620000 183.400000 146.820000 184.480000 ;
      RECT 58.620000 183.400000 101.820000 184.480000 ;
      RECT 13.620000 183.400000 56.820000 184.480000 ;
      RECT 7.860000 183.400000 11.820000 184.480000 ;
      RECT 0.000000 183.400000 5.260000 184.480000 ;
      RECT 0.000000 183.390000 548.960000 183.400000 ;
      RECT 0.000000 181.930000 550.160000 183.390000 ;
      RECT 0.000000 181.760000 548.960000 181.930000 ;
      RECT 547.900000 180.950000 548.960000 181.760000 ;
      RECT 547.900000 180.680000 550.160000 180.950000 ;
      RECT 506.620000 180.680000 545.300000 181.760000 ;
      RECT 461.620000 180.680000 504.820000 181.760000 ;
      RECT 416.620000 180.680000 459.820000 181.760000 ;
      RECT 371.620000 180.680000 414.820000 181.760000 ;
      RECT 326.620000 180.680000 369.820000 181.760000 ;
      RECT 281.620000 180.680000 324.820000 181.760000 ;
      RECT 236.620000 180.680000 279.820000 181.760000 ;
      RECT 191.620000 180.680000 234.820000 181.760000 ;
      RECT 146.620000 180.680000 189.820000 181.760000 ;
      RECT 101.620000 180.680000 144.820000 181.760000 ;
      RECT 56.620000 180.680000 99.820000 181.760000 ;
      RECT 11.620000 180.680000 54.820000 181.760000 ;
      RECT 4.860000 180.680000 9.655000 181.760000 ;
      RECT 0.000000 180.680000 2.260000 181.760000 ;
      RECT 0.000000 180.100000 550.160000 180.680000 ;
      RECT 0.000000 179.120000 548.960000 180.100000 ;
      RECT 0.000000 179.040000 550.160000 179.120000 ;
      RECT 544.900000 177.960000 550.160000 179.040000 ;
      RECT 508.620000 177.960000 542.300000 179.040000 ;
      RECT 463.620000 177.960000 506.820000 179.040000 ;
      RECT 418.620000 177.960000 461.820000 179.040000 ;
      RECT 373.620000 177.960000 416.820000 179.040000 ;
      RECT 328.620000 177.960000 371.820000 179.040000 ;
      RECT 283.620000 177.960000 326.820000 179.040000 ;
      RECT 238.620000 177.960000 281.820000 179.040000 ;
      RECT 193.620000 177.960000 236.820000 179.040000 ;
      RECT 148.620000 177.960000 191.820000 179.040000 ;
      RECT 103.620000 177.960000 146.820000 179.040000 ;
      RECT 58.620000 177.960000 101.820000 179.040000 ;
      RECT 13.620000 177.960000 56.820000 179.040000 ;
      RECT 7.860000 177.960000 11.820000 179.040000 ;
      RECT 0.000000 177.960000 5.260000 179.040000 ;
      RECT 0.000000 177.660000 550.160000 177.960000 ;
      RECT 0.000000 176.680000 548.960000 177.660000 ;
      RECT 0.000000 176.320000 550.160000 176.680000 ;
      RECT 547.900000 175.240000 550.160000 176.320000 ;
      RECT 506.620000 175.240000 545.300000 176.320000 ;
      RECT 461.620000 175.240000 504.820000 176.320000 ;
      RECT 416.620000 175.240000 459.820000 176.320000 ;
      RECT 371.620000 175.240000 414.820000 176.320000 ;
      RECT 326.620000 175.240000 369.820000 176.320000 ;
      RECT 281.620000 175.240000 324.820000 176.320000 ;
      RECT 236.620000 175.240000 279.820000 176.320000 ;
      RECT 191.620000 175.240000 234.820000 176.320000 ;
      RECT 146.620000 175.240000 189.820000 176.320000 ;
      RECT 101.620000 175.240000 144.820000 176.320000 ;
      RECT 56.620000 175.240000 99.820000 176.320000 ;
      RECT 11.620000 175.240000 54.820000 176.320000 ;
      RECT 4.860000 175.240000 9.655000 176.320000 ;
      RECT 0.000000 175.240000 2.260000 176.320000 ;
      RECT 0.000000 175.220000 550.160000 175.240000 ;
      RECT 0.000000 174.240000 548.960000 175.220000 ;
      RECT 0.000000 173.600000 550.160000 174.240000 ;
      RECT 544.900000 172.780000 550.160000 173.600000 ;
      RECT 544.900000 172.520000 548.960000 172.780000 ;
      RECT 508.620000 172.520000 542.300000 173.600000 ;
      RECT 463.620000 172.520000 506.820000 173.600000 ;
      RECT 418.620000 172.520000 461.820000 173.600000 ;
      RECT 373.620000 172.520000 416.820000 173.600000 ;
      RECT 328.620000 172.520000 371.820000 173.600000 ;
      RECT 283.620000 172.520000 326.820000 173.600000 ;
      RECT 238.620000 172.520000 281.820000 173.600000 ;
      RECT 193.620000 172.520000 236.820000 173.600000 ;
      RECT 148.620000 172.520000 191.820000 173.600000 ;
      RECT 103.620000 172.520000 146.820000 173.600000 ;
      RECT 58.620000 172.520000 101.820000 173.600000 ;
      RECT 13.620000 172.520000 56.820000 173.600000 ;
      RECT 7.860000 172.520000 11.820000 173.600000 ;
      RECT 0.000000 172.520000 5.260000 173.600000 ;
      RECT 0.000000 171.800000 548.960000 172.520000 ;
      RECT 0.000000 170.950000 550.160000 171.800000 ;
      RECT 0.000000 170.880000 548.960000 170.950000 ;
      RECT 547.900000 169.970000 548.960000 170.880000 ;
      RECT 547.900000 169.800000 550.160000 169.970000 ;
      RECT 506.620000 169.800000 545.300000 170.880000 ;
      RECT 461.620000 169.800000 504.820000 170.880000 ;
      RECT 416.620000 169.800000 459.820000 170.880000 ;
      RECT 371.620000 169.800000 414.820000 170.880000 ;
      RECT 326.620000 169.800000 369.820000 170.880000 ;
      RECT 281.620000 169.800000 324.820000 170.880000 ;
      RECT 236.620000 169.800000 279.820000 170.880000 ;
      RECT 191.620000 169.800000 234.820000 170.880000 ;
      RECT 146.620000 169.800000 189.820000 170.880000 ;
      RECT 101.620000 169.800000 144.820000 170.880000 ;
      RECT 56.620000 169.800000 99.820000 170.880000 ;
      RECT 11.620000 169.800000 54.820000 170.880000 ;
      RECT 4.860000 169.800000 9.655000 170.880000 ;
      RECT 0.000000 169.800000 2.260000 170.880000 ;
      RECT 0.000000 168.510000 550.160000 169.800000 ;
      RECT 0.000000 168.160000 548.960000 168.510000 ;
      RECT 544.900000 167.530000 548.960000 168.160000 ;
      RECT 544.900000 167.080000 550.160000 167.530000 ;
      RECT 508.620000 167.080000 542.300000 168.160000 ;
      RECT 463.620000 167.080000 506.820000 168.160000 ;
      RECT 418.620000 167.080000 461.820000 168.160000 ;
      RECT 373.620000 167.080000 416.820000 168.160000 ;
      RECT 328.620000 167.080000 371.820000 168.160000 ;
      RECT 283.620000 167.080000 326.820000 168.160000 ;
      RECT 238.620000 167.080000 281.820000 168.160000 ;
      RECT 193.620000 167.080000 236.820000 168.160000 ;
      RECT 148.620000 167.080000 191.820000 168.160000 ;
      RECT 103.620000 167.080000 146.820000 168.160000 ;
      RECT 58.620000 167.080000 101.820000 168.160000 ;
      RECT 13.620000 167.080000 56.820000 168.160000 ;
      RECT 7.860000 167.080000 11.820000 168.160000 ;
      RECT 0.000000 167.080000 5.260000 168.160000 ;
      RECT 0.000000 166.070000 550.160000 167.080000 ;
      RECT 0.000000 165.440000 548.960000 166.070000 ;
      RECT 547.900000 165.090000 548.960000 165.440000 ;
      RECT 547.900000 164.360000 550.160000 165.090000 ;
      RECT 506.620000 164.360000 545.300000 165.440000 ;
      RECT 461.620000 164.360000 504.820000 165.440000 ;
      RECT 416.620000 164.360000 459.820000 165.440000 ;
      RECT 371.620000 164.360000 414.820000 165.440000 ;
      RECT 326.620000 164.360000 369.820000 165.440000 ;
      RECT 281.620000 164.360000 324.820000 165.440000 ;
      RECT 236.620000 164.360000 279.820000 165.440000 ;
      RECT 191.620000 164.360000 234.820000 165.440000 ;
      RECT 146.620000 164.360000 189.820000 165.440000 ;
      RECT 101.620000 164.360000 144.820000 165.440000 ;
      RECT 56.620000 164.360000 99.820000 165.440000 ;
      RECT 11.620000 164.360000 54.820000 165.440000 ;
      RECT 4.860000 164.360000 9.655000 165.440000 ;
      RECT 0.000000 164.360000 2.260000 165.440000 ;
      RECT 0.000000 163.630000 550.160000 164.360000 ;
      RECT 0.000000 162.720000 548.960000 163.630000 ;
      RECT 544.900000 162.650000 548.960000 162.720000 ;
      RECT 544.900000 161.640000 550.160000 162.650000 ;
      RECT 508.620000 161.640000 542.300000 162.720000 ;
      RECT 463.620000 161.640000 506.820000 162.720000 ;
      RECT 418.620000 161.640000 461.820000 162.720000 ;
      RECT 373.620000 161.640000 416.820000 162.720000 ;
      RECT 328.620000 161.640000 371.820000 162.720000 ;
      RECT 283.620000 161.640000 326.820000 162.720000 ;
      RECT 238.620000 161.640000 281.820000 162.720000 ;
      RECT 193.620000 161.640000 236.820000 162.720000 ;
      RECT 148.620000 161.640000 191.820000 162.720000 ;
      RECT 103.620000 161.640000 146.820000 162.720000 ;
      RECT 58.620000 161.640000 101.820000 162.720000 ;
      RECT 13.620000 161.640000 56.820000 162.720000 ;
      RECT 7.860000 161.640000 11.820000 162.720000 ;
      RECT 0.000000 161.640000 5.260000 162.720000 ;
      RECT 0.000000 161.190000 550.160000 161.640000 ;
      RECT 0.000000 160.210000 548.960000 161.190000 ;
      RECT 0.000000 160.000000 550.160000 160.210000 ;
      RECT 547.900000 159.360000 550.160000 160.000000 ;
      RECT 547.900000 158.920000 548.960000 159.360000 ;
      RECT 506.620000 158.920000 545.300000 160.000000 ;
      RECT 461.620000 158.920000 504.820000 160.000000 ;
      RECT 416.620000 158.920000 459.820000 160.000000 ;
      RECT 371.620000 158.920000 414.820000 160.000000 ;
      RECT 326.620000 158.920000 369.820000 160.000000 ;
      RECT 281.620000 158.920000 324.820000 160.000000 ;
      RECT 236.620000 158.920000 279.820000 160.000000 ;
      RECT 191.620000 158.920000 234.820000 160.000000 ;
      RECT 146.620000 158.920000 189.820000 160.000000 ;
      RECT 101.620000 158.920000 144.820000 160.000000 ;
      RECT 56.620000 158.920000 99.820000 160.000000 ;
      RECT 11.620000 158.920000 54.820000 160.000000 ;
      RECT 4.860000 158.920000 9.655000 160.000000 ;
      RECT 0.000000 158.920000 2.260000 160.000000 ;
      RECT 0.000000 158.380000 548.960000 158.920000 ;
      RECT 0.000000 157.280000 550.160000 158.380000 ;
      RECT 544.900000 156.920000 550.160000 157.280000 ;
      RECT 544.900000 156.200000 548.960000 156.920000 ;
      RECT 508.620000 156.200000 542.300000 157.280000 ;
      RECT 463.620000 156.200000 506.820000 157.280000 ;
      RECT 418.620000 156.200000 461.820000 157.280000 ;
      RECT 373.620000 156.200000 416.820000 157.280000 ;
      RECT 328.620000 156.200000 371.820000 157.280000 ;
      RECT 283.620000 156.200000 326.820000 157.280000 ;
      RECT 238.620000 156.200000 281.820000 157.280000 ;
      RECT 193.620000 156.200000 236.820000 157.280000 ;
      RECT 148.620000 156.200000 191.820000 157.280000 ;
      RECT 103.620000 156.200000 146.820000 157.280000 ;
      RECT 58.620000 156.200000 101.820000 157.280000 ;
      RECT 13.620000 156.200000 56.820000 157.280000 ;
      RECT 7.860000 156.200000 11.820000 157.280000 ;
      RECT 0.000000 156.200000 5.260000 157.280000 ;
      RECT 0.000000 155.940000 548.960000 156.200000 ;
      RECT 0.000000 154.560000 550.160000 155.940000 ;
      RECT 547.900000 154.480000 550.160000 154.560000 ;
      RECT 547.900000 153.500000 548.960000 154.480000 ;
      RECT 547.900000 153.480000 550.160000 153.500000 ;
      RECT 506.620000 153.480000 545.300000 154.560000 ;
      RECT 461.620000 153.480000 504.820000 154.560000 ;
      RECT 416.620000 153.480000 459.820000 154.560000 ;
      RECT 371.620000 153.480000 414.820000 154.560000 ;
      RECT 326.620000 153.480000 369.820000 154.560000 ;
      RECT 281.620000 153.480000 324.820000 154.560000 ;
      RECT 236.620000 153.480000 279.820000 154.560000 ;
      RECT 191.620000 153.480000 234.820000 154.560000 ;
      RECT 146.620000 153.480000 189.820000 154.560000 ;
      RECT 101.620000 153.480000 144.820000 154.560000 ;
      RECT 56.620000 153.480000 99.820000 154.560000 ;
      RECT 11.620000 153.480000 54.820000 154.560000 ;
      RECT 4.860000 153.480000 9.655000 154.560000 ;
      RECT 0.000000 153.480000 2.260000 154.560000 ;
      RECT 0.000000 152.040000 550.160000 153.480000 ;
      RECT 0.000000 151.840000 548.960000 152.040000 ;
      RECT 544.900000 151.060000 548.960000 151.840000 ;
      RECT 544.900000 150.760000 550.160000 151.060000 ;
      RECT 508.620000 150.760000 542.300000 151.840000 ;
      RECT 463.620000 150.760000 506.820000 151.840000 ;
      RECT 418.620000 150.760000 461.820000 151.840000 ;
      RECT 373.620000 150.760000 416.820000 151.840000 ;
      RECT 328.620000 150.760000 371.820000 151.840000 ;
      RECT 283.620000 150.760000 326.820000 151.840000 ;
      RECT 238.620000 150.760000 281.820000 151.840000 ;
      RECT 193.620000 150.760000 236.820000 151.840000 ;
      RECT 148.620000 150.760000 191.820000 151.840000 ;
      RECT 103.620000 150.760000 146.820000 151.840000 ;
      RECT 58.620000 150.760000 101.820000 151.840000 ;
      RECT 13.620000 150.760000 56.820000 151.840000 ;
      RECT 7.860000 150.760000 11.820000 151.840000 ;
      RECT 0.000000 150.760000 5.260000 151.840000 ;
      RECT 0.000000 150.210000 550.160000 150.760000 ;
      RECT 0.000000 149.230000 548.960000 150.210000 ;
      RECT 0.000000 149.120000 550.160000 149.230000 ;
      RECT 547.900000 148.040000 550.160000 149.120000 ;
      RECT 506.620000 148.040000 545.300000 149.120000 ;
      RECT 461.620000 148.040000 504.820000 149.120000 ;
      RECT 416.620000 148.040000 459.820000 149.120000 ;
      RECT 371.620000 148.040000 414.820000 149.120000 ;
      RECT 326.620000 148.040000 369.820000 149.120000 ;
      RECT 281.620000 148.040000 324.820000 149.120000 ;
      RECT 236.620000 148.040000 279.820000 149.120000 ;
      RECT 191.620000 148.040000 234.820000 149.120000 ;
      RECT 146.620000 148.040000 189.820000 149.120000 ;
      RECT 101.620000 148.040000 144.820000 149.120000 ;
      RECT 56.620000 148.040000 99.820000 149.120000 ;
      RECT 11.620000 148.040000 54.820000 149.120000 ;
      RECT 4.860000 148.040000 9.655000 149.120000 ;
      RECT 0.000000 148.040000 2.260000 149.120000 ;
      RECT 0.000000 147.770000 550.160000 148.040000 ;
      RECT 0.000000 146.790000 548.960000 147.770000 ;
      RECT 0.000000 146.400000 550.160000 146.790000 ;
      RECT 544.900000 145.330000 550.160000 146.400000 ;
      RECT 544.900000 145.320000 548.960000 145.330000 ;
      RECT 508.620000 145.320000 542.300000 146.400000 ;
      RECT 463.620000 145.320000 506.820000 146.400000 ;
      RECT 418.620000 145.320000 461.820000 146.400000 ;
      RECT 373.620000 145.320000 416.820000 146.400000 ;
      RECT 328.620000 145.320000 371.820000 146.400000 ;
      RECT 283.620000 145.320000 326.820000 146.400000 ;
      RECT 238.620000 145.320000 281.820000 146.400000 ;
      RECT 193.620000 145.320000 236.820000 146.400000 ;
      RECT 148.620000 145.320000 191.820000 146.400000 ;
      RECT 103.620000 145.320000 146.820000 146.400000 ;
      RECT 58.620000 145.320000 101.820000 146.400000 ;
      RECT 13.620000 145.320000 56.820000 146.400000 ;
      RECT 7.860000 145.320000 11.820000 146.400000 ;
      RECT 0.000000 145.320000 5.260000 146.400000 ;
      RECT 0.000000 144.350000 548.960000 145.320000 ;
      RECT 0.000000 143.680000 550.160000 144.350000 ;
      RECT 547.900000 142.890000 550.160000 143.680000 ;
      RECT 547.900000 142.600000 548.960000 142.890000 ;
      RECT 506.620000 142.600000 545.300000 143.680000 ;
      RECT 461.620000 142.600000 504.820000 143.680000 ;
      RECT 416.620000 142.600000 459.820000 143.680000 ;
      RECT 371.620000 142.600000 414.820000 143.680000 ;
      RECT 326.620000 142.600000 369.820000 143.680000 ;
      RECT 281.620000 142.600000 324.820000 143.680000 ;
      RECT 236.620000 142.600000 279.820000 143.680000 ;
      RECT 191.620000 142.600000 234.820000 143.680000 ;
      RECT 146.620000 142.600000 189.820000 143.680000 ;
      RECT 101.620000 142.600000 144.820000 143.680000 ;
      RECT 56.620000 142.600000 99.820000 143.680000 ;
      RECT 11.620000 142.600000 54.820000 143.680000 ;
      RECT 4.860000 142.600000 9.655000 143.680000 ;
      RECT 0.000000 142.600000 2.260000 143.680000 ;
      RECT 0.000000 141.910000 548.960000 142.600000 ;
      RECT 0.000000 141.060000 550.160000 141.910000 ;
      RECT 0.000000 140.960000 548.960000 141.060000 ;
      RECT 544.900000 140.080000 548.960000 140.960000 ;
      RECT 544.900000 139.880000 550.160000 140.080000 ;
      RECT 508.620000 139.880000 542.300000 140.960000 ;
      RECT 463.620000 139.880000 506.820000 140.960000 ;
      RECT 418.620000 139.880000 461.820000 140.960000 ;
      RECT 373.620000 139.880000 416.820000 140.960000 ;
      RECT 328.620000 139.880000 371.820000 140.960000 ;
      RECT 283.620000 139.880000 326.820000 140.960000 ;
      RECT 238.620000 139.880000 281.820000 140.960000 ;
      RECT 193.620000 139.880000 236.820000 140.960000 ;
      RECT 148.620000 139.880000 191.820000 140.960000 ;
      RECT 103.620000 139.880000 146.820000 140.960000 ;
      RECT 58.620000 139.880000 101.820000 140.960000 ;
      RECT 13.620000 139.880000 56.820000 140.960000 ;
      RECT 7.860000 139.880000 11.820000 140.960000 ;
      RECT 0.000000 139.880000 5.260000 140.960000 ;
      RECT 0.000000 138.620000 550.160000 139.880000 ;
      RECT 0.000000 138.240000 548.960000 138.620000 ;
      RECT 547.900000 137.640000 548.960000 138.240000 ;
      RECT 547.900000 137.160000 550.160000 137.640000 ;
      RECT 506.620000 137.160000 545.300000 138.240000 ;
      RECT 461.620000 137.160000 504.820000 138.240000 ;
      RECT 416.620000 137.160000 459.820000 138.240000 ;
      RECT 371.620000 137.160000 414.820000 138.240000 ;
      RECT 326.620000 137.160000 369.820000 138.240000 ;
      RECT 281.620000 137.160000 324.820000 138.240000 ;
      RECT 236.620000 137.160000 279.820000 138.240000 ;
      RECT 191.620000 137.160000 234.820000 138.240000 ;
      RECT 146.620000 137.160000 189.820000 138.240000 ;
      RECT 101.620000 137.160000 144.820000 138.240000 ;
      RECT 56.620000 137.160000 99.820000 138.240000 ;
      RECT 11.620000 137.160000 54.820000 138.240000 ;
      RECT 4.860000 137.160000 9.655000 138.240000 ;
      RECT 0.000000 137.160000 2.260000 138.240000 ;
      RECT 0.000000 136.180000 550.160000 137.160000 ;
      RECT 0.000000 135.520000 548.960000 136.180000 ;
      RECT 544.900000 135.200000 548.960000 135.520000 ;
      RECT 544.900000 134.440000 550.160000 135.200000 ;
      RECT 508.620000 134.440000 542.300000 135.520000 ;
      RECT 463.620000 134.440000 506.820000 135.520000 ;
      RECT 418.620000 134.440000 461.820000 135.520000 ;
      RECT 373.620000 134.440000 416.820000 135.520000 ;
      RECT 328.620000 134.440000 371.820000 135.520000 ;
      RECT 283.620000 134.440000 326.820000 135.520000 ;
      RECT 238.620000 134.440000 281.820000 135.520000 ;
      RECT 193.620000 134.440000 236.820000 135.520000 ;
      RECT 148.620000 134.440000 191.820000 135.520000 ;
      RECT 103.620000 134.440000 146.820000 135.520000 ;
      RECT 58.620000 134.440000 101.820000 135.520000 ;
      RECT 13.620000 134.440000 56.820000 135.520000 ;
      RECT 7.860000 134.440000 11.820000 135.520000 ;
      RECT 0.000000 134.440000 5.260000 135.520000 ;
      RECT 0.000000 133.740000 550.160000 134.440000 ;
      RECT 0.000000 132.800000 548.960000 133.740000 ;
      RECT 547.900000 132.760000 548.960000 132.800000 ;
      RECT 547.900000 131.910000 550.160000 132.760000 ;
      RECT 547.900000 131.720000 548.960000 131.910000 ;
      RECT 506.620000 131.720000 545.300000 132.800000 ;
      RECT 461.620000 131.720000 504.820000 132.800000 ;
      RECT 416.620000 131.720000 459.820000 132.800000 ;
      RECT 371.620000 131.720000 414.820000 132.800000 ;
      RECT 326.620000 131.720000 369.820000 132.800000 ;
      RECT 281.620000 131.720000 324.820000 132.800000 ;
      RECT 236.620000 131.720000 279.820000 132.800000 ;
      RECT 191.620000 131.720000 234.820000 132.800000 ;
      RECT 146.620000 131.720000 189.820000 132.800000 ;
      RECT 101.620000 131.720000 144.820000 132.800000 ;
      RECT 56.620000 131.720000 99.820000 132.800000 ;
      RECT 11.620000 131.720000 54.820000 132.800000 ;
      RECT 4.860000 131.720000 9.655000 132.800000 ;
      RECT 0.000000 131.720000 2.260000 132.800000 ;
      RECT 0.000000 130.930000 548.960000 131.720000 ;
      RECT 0.000000 130.080000 550.160000 130.930000 ;
      RECT 544.900000 129.470000 550.160000 130.080000 ;
      RECT 544.900000 129.000000 548.960000 129.470000 ;
      RECT 508.620000 129.000000 542.300000 130.080000 ;
      RECT 463.620000 129.000000 506.820000 130.080000 ;
      RECT 418.620000 129.000000 461.820000 130.080000 ;
      RECT 373.620000 129.000000 416.820000 130.080000 ;
      RECT 328.620000 129.000000 371.820000 130.080000 ;
      RECT 283.620000 129.000000 326.820000 130.080000 ;
      RECT 238.620000 129.000000 281.820000 130.080000 ;
      RECT 193.620000 129.000000 236.820000 130.080000 ;
      RECT 148.620000 129.000000 191.820000 130.080000 ;
      RECT 103.620000 129.000000 146.820000 130.080000 ;
      RECT 58.620000 129.000000 101.820000 130.080000 ;
      RECT 13.620000 129.000000 56.820000 130.080000 ;
      RECT 7.860000 129.000000 11.820000 130.080000 ;
      RECT 0.000000 129.000000 5.260000 130.080000 ;
      RECT 0.000000 128.490000 548.960000 129.000000 ;
      RECT 0.000000 127.360000 550.160000 128.490000 ;
      RECT 547.900000 127.030000 550.160000 127.360000 ;
      RECT 547.900000 126.280000 548.960000 127.030000 ;
      RECT 506.620000 126.280000 545.300000 127.360000 ;
      RECT 461.620000 126.280000 504.820000 127.360000 ;
      RECT 416.620000 126.280000 459.820000 127.360000 ;
      RECT 371.620000 126.280000 414.820000 127.360000 ;
      RECT 326.620000 126.280000 369.820000 127.360000 ;
      RECT 281.620000 126.280000 324.820000 127.360000 ;
      RECT 236.620000 126.280000 279.820000 127.360000 ;
      RECT 191.620000 126.280000 234.820000 127.360000 ;
      RECT 146.620000 126.280000 189.820000 127.360000 ;
      RECT 101.620000 126.280000 144.820000 127.360000 ;
      RECT 56.620000 126.280000 99.820000 127.360000 ;
      RECT 11.620000 126.280000 54.820000 127.360000 ;
      RECT 4.860000 126.280000 9.655000 127.360000 ;
      RECT 0.000000 126.280000 2.260000 127.360000 ;
      RECT 0.000000 126.050000 548.960000 126.280000 ;
      RECT 0.000000 124.640000 550.160000 126.050000 ;
      RECT 544.900000 124.590000 550.160000 124.640000 ;
      RECT 544.900000 123.610000 548.960000 124.590000 ;
      RECT 544.900000 123.560000 550.160000 123.610000 ;
      RECT 508.620000 123.560000 542.300000 124.640000 ;
      RECT 463.620000 123.560000 506.820000 124.640000 ;
      RECT 418.620000 123.560000 461.820000 124.640000 ;
      RECT 373.620000 123.560000 416.820000 124.640000 ;
      RECT 328.620000 123.560000 371.820000 124.640000 ;
      RECT 283.620000 123.560000 326.820000 124.640000 ;
      RECT 238.620000 123.560000 281.820000 124.640000 ;
      RECT 193.620000 123.560000 236.820000 124.640000 ;
      RECT 148.620000 123.560000 191.820000 124.640000 ;
      RECT 103.620000 123.560000 146.820000 124.640000 ;
      RECT 58.620000 123.560000 101.820000 124.640000 ;
      RECT 13.620000 123.560000 56.820000 124.640000 ;
      RECT 7.860000 123.560000 11.820000 124.640000 ;
      RECT 0.000000 123.560000 5.260000 124.640000 ;
      RECT 0.000000 122.760000 550.160000 123.560000 ;
      RECT 0.000000 121.920000 548.960000 122.760000 ;
      RECT 547.900000 121.780000 548.960000 121.920000 ;
      RECT 547.900000 120.840000 550.160000 121.780000 ;
      RECT 506.620000 120.840000 545.300000 121.920000 ;
      RECT 461.620000 120.840000 504.820000 121.920000 ;
      RECT 416.620000 120.840000 459.820000 121.920000 ;
      RECT 371.620000 120.840000 414.820000 121.920000 ;
      RECT 326.620000 120.840000 369.820000 121.920000 ;
      RECT 281.620000 120.840000 324.820000 121.920000 ;
      RECT 236.620000 120.840000 279.820000 121.920000 ;
      RECT 191.620000 120.840000 234.820000 121.920000 ;
      RECT 146.620000 120.840000 189.820000 121.920000 ;
      RECT 101.620000 120.840000 144.820000 121.920000 ;
      RECT 56.620000 120.840000 99.820000 121.920000 ;
      RECT 11.620000 120.840000 54.820000 121.920000 ;
      RECT 4.860000 120.840000 9.655000 121.920000 ;
      RECT 0.000000 120.840000 2.260000 121.920000 ;
      RECT 0.000000 120.320000 550.160000 120.840000 ;
      RECT 0.000000 119.340000 548.960000 120.320000 ;
      RECT 0.000000 119.200000 550.160000 119.340000 ;
      RECT 544.900000 118.120000 550.160000 119.200000 ;
      RECT 508.620000 118.120000 542.300000 119.200000 ;
      RECT 463.620000 118.120000 506.820000 119.200000 ;
      RECT 418.620000 118.120000 461.820000 119.200000 ;
      RECT 373.620000 118.120000 416.820000 119.200000 ;
      RECT 328.620000 118.120000 371.820000 119.200000 ;
      RECT 283.620000 118.120000 326.820000 119.200000 ;
      RECT 238.620000 118.120000 281.820000 119.200000 ;
      RECT 193.620000 118.120000 236.820000 119.200000 ;
      RECT 148.620000 118.120000 191.820000 119.200000 ;
      RECT 103.620000 118.120000 146.820000 119.200000 ;
      RECT 58.620000 118.120000 101.820000 119.200000 ;
      RECT 13.620000 118.120000 56.820000 119.200000 ;
      RECT 7.860000 118.120000 11.820000 119.200000 ;
      RECT 0.000000 118.120000 5.260000 119.200000 ;
      RECT 0.000000 117.880000 550.160000 118.120000 ;
      RECT 0.000000 116.900000 548.960000 117.880000 ;
      RECT 0.000000 116.480000 550.160000 116.900000 ;
      RECT 547.900000 115.440000 550.160000 116.480000 ;
      RECT 547.900000 115.400000 548.960000 115.440000 ;
      RECT 506.620000 115.400000 545.300000 116.480000 ;
      RECT 461.620000 115.400000 504.820000 116.480000 ;
      RECT 416.620000 115.400000 459.820000 116.480000 ;
      RECT 371.620000 115.400000 414.820000 116.480000 ;
      RECT 326.620000 115.400000 369.820000 116.480000 ;
      RECT 281.620000 115.400000 324.820000 116.480000 ;
      RECT 236.620000 115.400000 279.820000 116.480000 ;
      RECT 191.620000 115.400000 234.820000 116.480000 ;
      RECT 146.620000 115.400000 189.820000 116.480000 ;
      RECT 101.620000 115.400000 144.820000 116.480000 ;
      RECT 56.620000 115.400000 99.820000 116.480000 ;
      RECT 11.620000 115.400000 54.820000 116.480000 ;
      RECT 4.860000 115.400000 9.655000 116.480000 ;
      RECT 0.000000 115.400000 2.260000 116.480000 ;
      RECT 0.000000 114.460000 548.960000 115.400000 ;
      RECT 0.000000 113.760000 550.160000 114.460000 ;
      RECT 544.900000 113.610000 550.160000 113.760000 ;
      RECT 544.900000 112.680000 548.960000 113.610000 ;
      RECT 508.620000 112.680000 542.300000 113.760000 ;
      RECT 463.620000 112.680000 506.820000 113.760000 ;
      RECT 418.620000 112.680000 461.820000 113.760000 ;
      RECT 373.620000 112.680000 416.820000 113.760000 ;
      RECT 328.620000 112.680000 371.820000 113.760000 ;
      RECT 283.620000 112.680000 326.820000 113.760000 ;
      RECT 238.620000 112.680000 281.820000 113.760000 ;
      RECT 193.620000 112.680000 236.820000 113.760000 ;
      RECT 148.620000 112.680000 191.820000 113.760000 ;
      RECT 103.620000 112.680000 146.820000 113.760000 ;
      RECT 58.620000 112.680000 101.820000 113.760000 ;
      RECT 13.620000 112.680000 56.820000 113.760000 ;
      RECT 7.860000 112.680000 11.820000 113.760000 ;
      RECT 0.000000 112.680000 5.260000 113.760000 ;
      RECT 0.000000 112.630000 548.960000 112.680000 ;
      RECT 0.000000 111.170000 550.160000 112.630000 ;
      RECT 0.000000 111.040000 548.960000 111.170000 ;
      RECT 547.900000 110.190000 548.960000 111.040000 ;
      RECT 547.900000 109.960000 550.160000 110.190000 ;
      RECT 506.620000 109.960000 545.300000 111.040000 ;
      RECT 461.620000 109.960000 504.820000 111.040000 ;
      RECT 416.620000 109.960000 459.820000 111.040000 ;
      RECT 371.620000 109.960000 414.820000 111.040000 ;
      RECT 326.620000 109.960000 369.820000 111.040000 ;
      RECT 281.620000 109.960000 324.820000 111.040000 ;
      RECT 236.620000 109.960000 279.820000 111.040000 ;
      RECT 191.620000 109.960000 234.820000 111.040000 ;
      RECT 146.620000 109.960000 189.820000 111.040000 ;
      RECT 101.620000 109.960000 144.820000 111.040000 ;
      RECT 56.620000 109.960000 99.820000 111.040000 ;
      RECT 11.620000 109.960000 54.820000 111.040000 ;
      RECT 4.860000 109.960000 9.655000 111.040000 ;
      RECT 0.000000 109.960000 2.260000 111.040000 ;
      RECT 0.000000 108.730000 550.160000 109.960000 ;
      RECT 0.000000 108.320000 548.960000 108.730000 ;
      RECT 544.900000 107.750000 548.960000 108.320000 ;
      RECT 544.900000 107.240000 550.160000 107.750000 ;
      RECT 508.620000 107.240000 542.300000 108.320000 ;
      RECT 463.620000 107.240000 506.820000 108.320000 ;
      RECT 418.620000 107.240000 461.820000 108.320000 ;
      RECT 373.620000 107.240000 416.820000 108.320000 ;
      RECT 328.620000 107.240000 371.820000 108.320000 ;
      RECT 283.620000 107.240000 326.820000 108.320000 ;
      RECT 238.620000 107.240000 281.820000 108.320000 ;
      RECT 193.620000 107.240000 236.820000 108.320000 ;
      RECT 148.620000 107.240000 191.820000 108.320000 ;
      RECT 103.620000 107.240000 146.820000 108.320000 ;
      RECT 58.620000 107.240000 101.820000 108.320000 ;
      RECT 13.620000 107.240000 56.820000 108.320000 ;
      RECT 7.860000 107.240000 11.820000 108.320000 ;
      RECT 0.000000 107.240000 5.260000 108.320000 ;
      RECT 0.000000 106.290000 550.160000 107.240000 ;
      RECT 0.000000 105.600000 548.960000 106.290000 ;
      RECT 547.900000 105.310000 548.960000 105.600000 ;
      RECT 547.900000 104.520000 550.160000 105.310000 ;
      RECT 506.620000 104.520000 545.300000 105.600000 ;
      RECT 461.620000 104.520000 504.820000 105.600000 ;
      RECT 416.620000 104.520000 459.820000 105.600000 ;
      RECT 371.620000 104.520000 414.820000 105.600000 ;
      RECT 326.620000 104.520000 369.820000 105.600000 ;
      RECT 281.620000 104.520000 324.820000 105.600000 ;
      RECT 236.620000 104.520000 279.820000 105.600000 ;
      RECT 191.620000 104.520000 234.820000 105.600000 ;
      RECT 146.620000 104.520000 189.820000 105.600000 ;
      RECT 101.620000 104.520000 144.820000 105.600000 ;
      RECT 56.620000 104.520000 99.820000 105.600000 ;
      RECT 11.620000 104.520000 54.820000 105.600000 ;
      RECT 4.860000 104.520000 9.655000 105.600000 ;
      RECT 0.000000 104.520000 2.260000 105.600000 ;
      RECT 0.000000 104.460000 550.160000 104.520000 ;
      RECT 0.000000 103.480000 548.960000 104.460000 ;
      RECT 0.000000 102.880000 550.160000 103.480000 ;
      RECT 544.900000 102.020000 550.160000 102.880000 ;
      RECT 544.900000 101.800000 548.960000 102.020000 ;
      RECT 508.620000 101.800000 542.300000 102.880000 ;
      RECT 463.620000 101.800000 506.820000 102.880000 ;
      RECT 418.620000 101.800000 461.820000 102.880000 ;
      RECT 373.620000 101.800000 416.820000 102.880000 ;
      RECT 328.620000 101.800000 371.820000 102.880000 ;
      RECT 283.620000 101.800000 326.820000 102.880000 ;
      RECT 238.620000 101.800000 281.820000 102.880000 ;
      RECT 193.620000 101.800000 236.820000 102.880000 ;
      RECT 148.620000 101.800000 191.820000 102.880000 ;
      RECT 103.620000 101.800000 146.820000 102.880000 ;
      RECT 58.620000 101.800000 101.820000 102.880000 ;
      RECT 13.620000 101.800000 56.820000 102.880000 ;
      RECT 7.860000 101.800000 11.820000 102.880000 ;
      RECT 0.000000 101.800000 5.260000 102.880000 ;
      RECT 0.000000 101.040000 548.960000 101.800000 ;
      RECT 0.000000 100.160000 550.160000 101.040000 ;
      RECT 547.900000 99.580000 550.160000 100.160000 ;
      RECT 547.900000 99.080000 548.960000 99.580000 ;
      RECT 506.620000 99.080000 545.300000 100.160000 ;
      RECT 461.620000 99.080000 504.820000 100.160000 ;
      RECT 416.620000 99.080000 459.820000 100.160000 ;
      RECT 371.620000 99.080000 414.820000 100.160000 ;
      RECT 326.620000 99.080000 369.820000 100.160000 ;
      RECT 281.620000 99.080000 324.820000 100.160000 ;
      RECT 236.620000 99.080000 279.820000 100.160000 ;
      RECT 191.620000 99.080000 234.820000 100.160000 ;
      RECT 146.620000 99.080000 189.820000 100.160000 ;
      RECT 101.620000 99.080000 144.820000 100.160000 ;
      RECT 56.620000 99.080000 99.820000 100.160000 ;
      RECT 11.620000 99.080000 54.820000 100.160000 ;
      RECT 4.860000 99.080000 9.655000 100.160000 ;
      RECT 0.000000 99.080000 2.260000 100.160000 ;
      RECT 0.000000 98.600000 548.960000 99.080000 ;
      RECT 0.000000 97.440000 550.160000 98.600000 ;
      RECT 544.900000 97.140000 550.160000 97.440000 ;
      RECT 544.900000 96.360000 548.960000 97.140000 ;
      RECT 508.620000 96.360000 542.300000 97.440000 ;
      RECT 463.620000 96.360000 506.820000 97.440000 ;
      RECT 418.620000 96.360000 461.820000 97.440000 ;
      RECT 373.620000 96.360000 416.820000 97.440000 ;
      RECT 328.620000 96.360000 371.820000 97.440000 ;
      RECT 283.620000 96.360000 326.820000 97.440000 ;
      RECT 238.620000 96.360000 281.820000 97.440000 ;
      RECT 193.620000 96.360000 236.820000 97.440000 ;
      RECT 148.620000 96.360000 191.820000 97.440000 ;
      RECT 103.620000 96.360000 146.820000 97.440000 ;
      RECT 58.620000 96.360000 101.820000 97.440000 ;
      RECT 13.620000 96.360000 56.820000 97.440000 ;
      RECT 7.860000 96.360000 11.820000 97.440000 ;
      RECT 0.000000 96.360000 5.260000 97.440000 ;
      RECT 0.000000 96.160000 548.960000 96.360000 ;
      RECT 0.000000 95.310000 550.160000 96.160000 ;
      RECT 0.000000 94.720000 548.960000 95.310000 ;
      RECT 547.900000 94.330000 548.960000 94.720000 ;
      RECT 547.900000 93.640000 550.160000 94.330000 ;
      RECT 506.620000 93.640000 545.300000 94.720000 ;
      RECT 461.620000 93.640000 504.820000 94.720000 ;
      RECT 416.620000 93.640000 459.820000 94.720000 ;
      RECT 371.620000 93.640000 414.820000 94.720000 ;
      RECT 326.620000 93.640000 369.820000 94.720000 ;
      RECT 281.620000 93.640000 324.820000 94.720000 ;
      RECT 236.620000 93.640000 279.820000 94.720000 ;
      RECT 191.620000 93.640000 234.820000 94.720000 ;
      RECT 146.620000 93.640000 189.820000 94.720000 ;
      RECT 101.620000 93.640000 144.820000 94.720000 ;
      RECT 56.620000 93.640000 99.820000 94.720000 ;
      RECT 11.620000 93.640000 54.820000 94.720000 ;
      RECT 4.860000 93.640000 9.655000 94.720000 ;
      RECT 0.000000 93.640000 2.260000 94.720000 ;
      RECT 0.000000 92.870000 550.160000 93.640000 ;
      RECT 0.000000 92.000000 548.960000 92.870000 ;
      RECT 544.900000 91.890000 548.960000 92.000000 ;
      RECT 544.900000 90.920000 550.160000 91.890000 ;
      RECT 508.620000 90.920000 542.300000 92.000000 ;
      RECT 463.620000 90.920000 506.820000 92.000000 ;
      RECT 418.620000 90.920000 461.820000 92.000000 ;
      RECT 373.620000 90.920000 416.820000 92.000000 ;
      RECT 328.620000 90.920000 371.820000 92.000000 ;
      RECT 283.620000 90.920000 326.820000 92.000000 ;
      RECT 238.620000 90.920000 281.820000 92.000000 ;
      RECT 193.620000 90.920000 236.820000 92.000000 ;
      RECT 148.620000 90.920000 191.820000 92.000000 ;
      RECT 103.620000 90.920000 146.820000 92.000000 ;
      RECT 58.620000 90.920000 101.820000 92.000000 ;
      RECT 13.620000 90.920000 56.820000 92.000000 ;
      RECT 7.860000 90.920000 11.820000 92.000000 ;
      RECT 0.000000 90.920000 5.260000 92.000000 ;
      RECT 0.000000 90.430000 550.160000 90.920000 ;
      RECT 0.000000 89.450000 548.960000 90.430000 ;
      RECT 0.000000 89.280000 550.160000 89.450000 ;
      RECT 547.900000 88.200000 550.160000 89.280000 ;
      RECT 506.620000 88.200000 545.300000 89.280000 ;
      RECT 461.620000 88.200000 504.820000 89.280000 ;
      RECT 416.620000 88.200000 459.820000 89.280000 ;
      RECT 371.620000 88.200000 414.820000 89.280000 ;
      RECT 326.620000 88.200000 369.820000 89.280000 ;
      RECT 281.620000 88.200000 324.820000 89.280000 ;
      RECT 236.620000 88.200000 279.820000 89.280000 ;
      RECT 191.620000 88.200000 234.820000 89.280000 ;
      RECT 146.620000 88.200000 189.820000 89.280000 ;
      RECT 101.620000 88.200000 144.820000 89.280000 ;
      RECT 56.620000 88.200000 99.820000 89.280000 ;
      RECT 11.620000 88.200000 54.820000 89.280000 ;
      RECT 4.860000 88.200000 9.655000 89.280000 ;
      RECT 0.000000 88.200000 2.260000 89.280000 ;
      RECT 0.000000 87.990000 550.160000 88.200000 ;
      RECT 0.000000 87.010000 548.960000 87.990000 ;
      RECT 0.000000 86.560000 550.160000 87.010000 ;
      RECT 544.900000 85.550000 550.160000 86.560000 ;
      RECT 544.900000 85.480000 548.960000 85.550000 ;
      RECT 508.620000 85.480000 542.300000 86.560000 ;
      RECT 463.620000 85.480000 506.820000 86.560000 ;
      RECT 418.620000 85.480000 461.820000 86.560000 ;
      RECT 373.620000 85.480000 416.820000 86.560000 ;
      RECT 328.620000 85.480000 371.820000 86.560000 ;
      RECT 283.620000 85.480000 326.820000 86.560000 ;
      RECT 238.620000 85.480000 281.820000 86.560000 ;
      RECT 193.620000 85.480000 236.820000 86.560000 ;
      RECT 148.620000 85.480000 191.820000 86.560000 ;
      RECT 103.620000 85.480000 146.820000 86.560000 ;
      RECT 58.620000 85.480000 101.820000 86.560000 ;
      RECT 13.620000 85.480000 56.820000 86.560000 ;
      RECT 7.860000 85.480000 11.820000 86.560000 ;
      RECT 0.000000 85.480000 5.260000 86.560000 ;
      RECT 0.000000 84.570000 548.960000 85.480000 ;
      RECT 0.000000 83.840000 550.160000 84.570000 ;
      RECT 547.900000 83.720000 550.160000 83.840000 ;
      RECT 547.900000 82.760000 548.960000 83.720000 ;
      RECT 506.620000 82.760000 545.300000 83.840000 ;
      RECT 461.620000 82.760000 504.820000 83.840000 ;
      RECT 416.620000 82.760000 459.820000 83.840000 ;
      RECT 371.620000 82.760000 414.820000 83.840000 ;
      RECT 326.620000 82.760000 369.820000 83.840000 ;
      RECT 281.620000 82.760000 324.820000 83.840000 ;
      RECT 236.620000 82.760000 279.820000 83.840000 ;
      RECT 191.620000 82.760000 234.820000 83.840000 ;
      RECT 146.620000 82.760000 189.820000 83.840000 ;
      RECT 101.620000 82.760000 144.820000 83.840000 ;
      RECT 56.620000 82.760000 99.820000 83.840000 ;
      RECT 11.620000 82.760000 54.820000 83.840000 ;
      RECT 4.860000 82.760000 9.655000 83.840000 ;
      RECT 0.000000 82.760000 2.260000 83.840000 ;
      RECT 0.000000 82.740000 548.960000 82.760000 ;
      RECT 0.000000 81.280000 550.160000 82.740000 ;
      RECT 0.000000 81.120000 548.960000 81.280000 ;
      RECT 544.900000 80.300000 548.960000 81.120000 ;
      RECT 544.900000 80.040000 550.160000 80.300000 ;
      RECT 508.620000 80.040000 542.300000 81.120000 ;
      RECT 463.620000 80.040000 506.820000 81.120000 ;
      RECT 418.620000 80.040000 461.820000 81.120000 ;
      RECT 373.620000 80.040000 416.820000 81.120000 ;
      RECT 328.620000 80.040000 371.820000 81.120000 ;
      RECT 283.620000 80.040000 326.820000 81.120000 ;
      RECT 238.620000 80.040000 281.820000 81.120000 ;
      RECT 193.620000 80.040000 236.820000 81.120000 ;
      RECT 148.620000 80.040000 191.820000 81.120000 ;
      RECT 103.620000 80.040000 146.820000 81.120000 ;
      RECT 58.620000 80.040000 101.820000 81.120000 ;
      RECT 13.620000 80.040000 56.820000 81.120000 ;
      RECT 7.860000 80.040000 11.820000 81.120000 ;
      RECT 0.000000 80.040000 5.260000 81.120000 ;
      RECT 0.000000 78.840000 550.160000 80.040000 ;
      RECT 0.000000 78.400000 548.960000 78.840000 ;
      RECT 547.900000 77.860000 548.960000 78.400000 ;
      RECT 547.900000 77.320000 550.160000 77.860000 ;
      RECT 506.620000 77.320000 545.300000 78.400000 ;
      RECT 461.620000 77.320000 504.820000 78.400000 ;
      RECT 416.620000 77.320000 459.820000 78.400000 ;
      RECT 371.620000 77.320000 414.820000 78.400000 ;
      RECT 326.620000 77.320000 369.820000 78.400000 ;
      RECT 281.620000 77.320000 324.820000 78.400000 ;
      RECT 236.620000 77.320000 279.820000 78.400000 ;
      RECT 191.620000 77.320000 234.820000 78.400000 ;
      RECT 146.620000 77.320000 189.820000 78.400000 ;
      RECT 101.620000 77.320000 144.820000 78.400000 ;
      RECT 56.620000 77.320000 99.820000 78.400000 ;
      RECT 11.620000 77.320000 54.820000 78.400000 ;
      RECT 4.860000 77.320000 9.655000 78.400000 ;
      RECT 0.000000 77.320000 2.260000 78.400000 ;
      RECT 0.000000 76.400000 550.160000 77.320000 ;
      RECT 0.000000 75.680000 548.960000 76.400000 ;
      RECT 544.900000 75.420000 548.960000 75.680000 ;
      RECT 544.900000 74.600000 550.160000 75.420000 ;
      RECT 508.620000 74.600000 542.300000 75.680000 ;
      RECT 463.620000 74.600000 506.820000 75.680000 ;
      RECT 418.620000 74.600000 461.820000 75.680000 ;
      RECT 373.620000 74.600000 416.820000 75.680000 ;
      RECT 328.620000 74.600000 371.820000 75.680000 ;
      RECT 283.620000 74.600000 326.820000 75.680000 ;
      RECT 238.620000 74.600000 281.820000 75.680000 ;
      RECT 193.620000 74.600000 236.820000 75.680000 ;
      RECT 148.620000 74.600000 191.820000 75.680000 ;
      RECT 103.620000 74.600000 146.820000 75.680000 ;
      RECT 58.620000 74.600000 101.820000 75.680000 ;
      RECT 13.620000 74.600000 56.820000 75.680000 ;
      RECT 7.860000 74.600000 11.820000 75.680000 ;
      RECT 0.000000 74.600000 5.260000 75.680000 ;
      RECT 0.000000 74.570000 550.160000 74.600000 ;
      RECT 0.000000 73.590000 548.960000 74.570000 ;
      RECT 0.000000 72.960000 550.160000 73.590000 ;
      RECT 547.900000 72.130000 550.160000 72.960000 ;
      RECT 547.900000 71.880000 548.960000 72.130000 ;
      RECT 506.620000 71.880000 545.300000 72.960000 ;
      RECT 461.620000 71.880000 504.820000 72.960000 ;
      RECT 416.620000 71.880000 459.820000 72.960000 ;
      RECT 371.620000 71.880000 414.820000 72.960000 ;
      RECT 326.620000 71.880000 369.820000 72.960000 ;
      RECT 281.620000 71.880000 324.820000 72.960000 ;
      RECT 236.620000 71.880000 279.820000 72.960000 ;
      RECT 191.620000 71.880000 234.820000 72.960000 ;
      RECT 146.620000 71.880000 189.820000 72.960000 ;
      RECT 101.620000 71.880000 144.820000 72.960000 ;
      RECT 56.620000 71.880000 99.820000 72.960000 ;
      RECT 11.620000 71.880000 54.820000 72.960000 ;
      RECT 4.860000 71.880000 9.655000 72.960000 ;
      RECT 0.000000 71.880000 2.260000 72.960000 ;
      RECT 0.000000 71.150000 548.960000 71.880000 ;
      RECT 0.000000 70.240000 550.160000 71.150000 ;
      RECT 544.900000 69.690000 550.160000 70.240000 ;
      RECT 544.900000 69.160000 548.960000 69.690000 ;
      RECT 508.620000 69.160000 542.300000 70.240000 ;
      RECT 463.620000 69.160000 506.820000 70.240000 ;
      RECT 418.620000 69.160000 461.820000 70.240000 ;
      RECT 373.620000 69.160000 416.820000 70.240000 ;
      RECT 328.620000 69.160000 371.820000 70.240000 ;
      RECT 283.620000 69.160000 326.820000 70.240000 ;
      RECT 238.620000 69.160000 281.820000 70.240000 ;
      RECT 193.620000 69.160000 236.820000 70.240000 ;
      RECT 148.620000 69.160000 191.820000 70.240000 ;
      RECT 103.620000 69.160000 146.820000 70.240000 ;
      RECT 58.620000 69.160000 101.820000 70.240000 ;
      RECT 13.620000 69.160000 56.820000 70.240000 ;
      RECT 7.860000 69.160000 11.820000 70.240000 ;
      RECT 0.000000 69.160000 5.260000 70.240000 ;
      RECT 0.000000 68.710000 548.960000 69.160000 ;
      RECT 0.000000 67.520000 550.160000 68.710000 ;
      RECT 547.900000 67.250000 550.160000 67.520000 ;
      RECT 547.900000 66.440000 548.960000 67.250000 ;
      RECT 506.620000 66.440000 545.300000 67.520000 ;
      RECT 461.620000 66.440000 504.820000 67.520000 ;
      RECT 416.620000 66.440000 459.820000 67.520000 ;
      RECT 371.620000 66.440000 414.820000 67.520000 ;
      RECT 326.620000 66.440000 369.820000 67.520000 ;
      RECT 281.620000 66.440000 324.820000 67.520000 ;
      RECT 236.620000 66.440000 279.820000 67.520000 ;
      RECT 191.620000 66.440000 234.820000 67.520000 ;
      RECT 146.620000 66.440000 189.820000 67.520000 ;
      RECT 101.620000 66.440000 144.820000 67.520000 ;
      RECT 56.620000 66.440000 99.820000 67.520000 ;
      RECT 11.620000 66.440000 54.820000 67.520000 ;
      RECT 4.860000 66.440000 9.655000 67.520000 ;
      RECT 0.000000 66.440000 2.260000 67.520000 ;
      RECT 0.000000 66.270000 548.960000 66.440000 ;
      RECT 0.000000 65.420000 550.160000 66.270000 ;
      RECT 0.000000 64.800000 548.960000 65.420000 ;
      RECT 544.900000 64.440000 548.960000 64.800000 ;
      RECT 544.900000 63.720000 550.160000 64.440000 ;
      RECT 508.620000 63.720000 542.300000 64.800000 ;
      RECT 463.620000 63.720000 506.820000 64.800000 ;
      RECT 418.620000 63.720000 461.820000 64.800000 ;
      RECT 373.620000 63.720000 416.820000 64.800000 ;
      RECT 328.620000 63.720000 371.820000 64.800000 ;
      RECT 283.620000 63.720000 326.820000 64.800000 ;
      RECT 238.620000 63.720000 281.820000 64.800000 ;
      RECT 193.620000 63.720000 236.820000 64.800000 ;
      RECT 148.620000 63.720000 191.820000 64.800000 ;
      RECT 103.620000 63.720000 146.820000 64.800000 ;
      RECT 58.620000 63.720000 101.820000 64.800000 ;
      RECT 13.620000 63.720000 56.820000 64.800000 ;
      RECT 7.860000 63.720000 11.820000 64.800000 ;
      RECT 0.000000 63.720000 5.260000 64.800000 ;
      RECT 0.000000 62.980000 550.160000 63.720000 ;
      RECT 0.000000 62.080000 548.960000 62.980000 ;
      RECT 547.900000 62.000000 548.960000 62.080000 ;
      RECT 547.900000 61.000000 550.160000 62.000000 ;
      RECT 506.620000 61.000000 545.300000 62.080000 ;
      RECT 461.620000 61.000000 504.820000 62.080000 ;
      RECT 416.620000 61.000000 459.820000 62.080000 ;
      RECT 371.620000 61.000000 414.820000 62.080000 ;
      RECT 326.620000 61.000000 369.820000 62.080000 ;
      RECT 281.620000 61.000000 324.820000 62.080000 ;
      RECT 236.620000 61.000000 279.820000 62.080000 ;
      RECT 191.620000 61.000000 234.820000 62.080000 ;
      RECT 146.620000 61.000000 189.820000 62.080000 ;
      RECT 101.620000 61.000000 144.820000 62.080000 ;
      RECT 56.620000 61.000000 99.820000 62.080000 ;
      RECT 11.620000 61.000000 54.820000 62.080000 ;
      RECT 4.860000 61.000000 9.655000 62.080000 ;
      RECT 0.000000 61.000000 2.260000 62.080000 ;
      RECT 0.000000 60.540000 550.160000 61.000000 ;
      RECT 0.000000 59.560000 548.960000 60.540000 ;
      RECT 0.000000 59.360000 550.160000 59.560000 ;
      RECT 544.900000 58.280000 550.160000 59.360000 ;
      RECT 508.620000 58.280000 542.300000 59.360000 ;
      RECT 463.620000 58.280000 506.820000 59.360000 ;
      RECT 418.620000 58.280000 461.820000 59.360000 ;
      RECT 373.620000 58.280000 416.820000 59.360000 ;
      RECT 328.620000 58.280000 371.820000 59.360000 ;
      RECT 283.620000 58.280000 326.820000 59.360000 ;
      RECT 238.620000 58.280000 281.820000 59.360000 ;
      RECT 193.620000 58.280000 236.820000 59.360000 ;
      RECT 148.620000 58.280000 191.820000 59.360000 ;
      RECT 103.620000 58.280000 146.820000 59.360000 ;
      RECT 58.620000 58.280000 101.820000 59.360000 ;
      RECT 13.620000 58.280000 56.820000 59.360000 ;
      RECT 7.860000 58.280000 11.820000 59.360000 ;
      RECT 0.000000 58.280000 5.260000 59.360000 ;
      RECT 0.000000 58.100000 550.160000 58.280000 ;
      RECT 0.000000 57.120000 548.960000 58.100000 ;
      RECT 0.000000 56.640000 550.160000 57.120000 ;
      RECT 547.900000 56.270000 550.160000 56.640000 ;
      RECT 547.900000 55.560000 548.960000 56.270000 ;
      RECT 506.620000 55.560000 545.300000 56.640000 ;
      RECT 461.620000 55.560000 504.820000 56.640000 ;
      RECT 416.620000 55.560000 459.820000 56.640000 ;
      RECT 371.620000 55.560000 414.820000 56.640000 ;
      RECT 326.620000 55.560000 369.820000 56.640000 ;
      RECT 281.620000 55.560000 324.820000 56.640000 ;
      RECT 236.620000 55.560000 279.820000 56.640000 ;
      RECT 191.620000 55.560000 234.820000 56.640000 ;
      RECT 146.620000 55.560000 189.820000 56.640000 ;
      RECT 101.620000 55.560000 144.820000 56.640000 ;
      RECT 56.620000 55.560000 99.820000 56.640000 ;
      RECT 11.620000 55.560000 54.820000 56.640000 ;
      RECT 4.860000 55.560000 9.655000 56.640000 ;
      RECT 0.000000 55.560000 2.260000 56.640000 ;
      RECT 0.000000 55.290000 548.960000 55.560000 ;
      RECT 0.000000 53.920000 550.160000 55.290000 ;
      RECT 544.900000 53.830000 550.160000 53.920000 ;
      RECT 544.900000 52.850000 548.960000 53.830000 ;
      RECT 544.900000 52.840000 550.160000 52.850000 ;
      RECT 508.620000 52.840000 542.300000 53.920000 ;
      RECT 463.620000 52.840000 506.820000 53.920000 ;
      RECT 418.620000 52.840000 461.820000 53.920000 ;
      RECT 373.620000 52.840000 416.820000 53.920000 ;
      RECT 328.620000 52.840000 371.820000 53.920000 ;
      RECT 283.620000 52.840000 326.820000 53.920000 ;
      RECT 238.620000 52.840000 281.820000 53.920000 ;
      RECT 193.620000 52.840000 236.820000 53.920000 ;
      RECT 148.620000 52.840000 191.820000 53.920000 ;
      RECT 103.620000 52.840000 146.820000 53.920000 ;
      RECT 58.620000 52.840000 101.820000 53.920000 ;
      RECT 13.620000 52.840000 56.820000 53.920000 ;
      RECT 7.860000 52.840000 11.820000 53.920000 ;
      RECT 0.000000 52.840000 5.260000 53.920000 ;
      RECT 0.000000 51.390000 550.160000 52.840000 ;
      RECT 0.000000 51.200000 548.960000 51.390000 ;
      RECT 547.900000 50.410000 548.960000 51.200000 ;
      RECT 547.900000 50.120000 550.160000 50.410000 ;
      RECT 506.620000 50.120000 545.300000 51.200000 ;
      RECT 461.620000 50.120000 504.820000 51.200000 ;
      RECT 416.620000 50.120000 459.820000 51.200000 ;
      RECT 371.620000 50.120000 414.820000 51.200000 ;
      RECT 326.620000 50.120000 369.820000 51.200000 ;
      RECT 281.620000 50.120000 324.820000 51.200000 ;
      RECT 236.620000 50.120000 279.820000 51.200000 ;
      RECT 191.620000 50.120000 234.820000 51.200000 ;
      RECT 146.620000 50.120000 189.820000 51.200000 ;
      RECT 101.620000 50.120000 144.820000 51.200000 ;
      RECT 56.620000 50.120000 99.820000 51.200000 ;
      RECT 11.620000 50.120000 54.820000 51.200000 ;
      RECT 4.860000 50.120000 9.655000 51.200000 ;
      RECT 0.000000 50.120000 2.260000 51.200000 ;
      RECT 0.000000 48.950000 550.160000 50.120000 ;
      RECT 0.000000 48.480000 548.960000 48.950000 ;
      RECT 544.900000 47.970000 548.960000 48.480000 ;
      RECT 544.900000 47.400000 550.160000 47.970000 ;
      RECT 508.620000 47.400000 542.300000 48.480000 ;
      RECT 463.620000 47.400000 506.820000 48.480000 ;
      RECT 418.620000 47.400000 461.820000 48.480000 ;
      RECT 373.620000 47.400000 416.820000 48.480000 ;
      RECT 328.620000 47.400000 371.820000 48.480000 ;
      RECT 283.620000 47.400000 326.820000 48.480000 ;
      RECT 238.620000 47.400000 281.820000 48.480000 ;
      RECT 193.620000 47.400000 236.820000 48.480000 ;
      RECT 148.620000 47.400000 191.820000 48.480000 ;
      RECT 103.620000 47.400000 146.820000 48.480000 ;
      RECT 58.620000 47.400000 101.820000 48.480000 ;
      RECT 13.620000 47.400000 56.820000 48.480000 ;
      RECT 7.860000 47.400000 11.820000 48.480000 ;
      RECT 0.000000 47.400000 5.260000 48.480000 ;
      RECT 0.000000 47.120000 550.160000 47.400000 ;
      RECT 0.000000 46.140000 548.960000 47.120000 ;
      RECT 0.000000 45.760000 550.160000 46.140000 ;
      RECT 547.900000 44.680000 550.160000 45.760000 ;
      RECT 506.620000 44.680000 545.300000 45.760000 ;
      RECT 461.620000 44.680000 504.820000 45.760000 ;
      RECT 416.620000 44.680000 459.820000 45.760000 ;
      RECT 371.620000 44.680000 414.820000 45.760000 ;
      RECT 326.620000 44.680000 369.820000 45.760000 ;
      RECT 281.620000 44.680000 324.820000 45.760000 ;
      RECT 236.620000 44.680000 279.820000 45.760000 ;
      RECT 191.620000 44.680000 234.820000 45.760000 ;
      RECT 146.620000 44.680000 189.820000 45.760000 ;
      RECT 101.620000 44.680000 144.820000 45.760000 ;
      RECT 56.620000 44.680000 99.820000 45.760000 ;
      RECT 11.620000 44.680000 54.820000 45.760000 ;
      RECT 4.860000 44.680000 9.655000 45.760000 ;
      RECT 0.000000 44.680000 2.260000 45.760000 ;
      RECT 0.000000 43.700000 548.960000 44.680000 ;
      RECT 0.000000 43.040000 550.160000 43.700000 ;
      RECT 544.900000 42.240000 550.160000 43.040000 ;
      RECT 544.900000 41.960000 548.960000 42.240000 ;
      RECT 508.620000 41.960000 542.300000 43.040000 ;
      RECT 463.620000 41.960000 506.820000 43.040000 ;
      RECT 418.620000 41.960000 461.820000 43.040000 ;
      RECT 373.620000 41.960000 416.820000 43.040000 ;
      RECT 328.620000 41.960000 371.820000 43.040000 ;
      RECT 283.620000 41.960000 326.820000 43.040000 ;
      RECT 238.620000 41.960000 281.820000 43.040000 ;
      RECT 193.620000 41.960000 236.820000 43.040000 ;
      RECT 148.620000 41.960000 191.820000 43.040000 ;
      RECT 103.620000 41.960000 146.820000 43.040000 ;
      RECT 58.620000 41.960000 101.820000 43.040000 ;
      RECT 13.620000 41.960000 56.820000 43.040000 ;
      RECT 7.860000 41.960000 11.820000 43.040000 ;
      RECT 0.000000 41.960000 5.260000 43.040000 ;
      RECT 0.000000 41.260000 548.960000 41.960000 ;
      RECT 0.000000 40.320000 550.160000 41.260000 ;
      RECT 547.900000 39.800000 550.160000 40.320000 ;
      RECT 547.900000 39.240000 548.960000 39.800000 ;
      RECT 506.620000 39.240000 545.300000 40.320000 ;
      RECT 461.620000 39.240000 504.820000 40.320000 ;
      RECT 416.620000 39.240000 459.820000 40.320000 ;
      RECT 371.620000 39.240000 414.820000 40.320000 ;
      RECT 326.620000 39.240000 369.820000 40.320000 ;
      RECT 281.620000 39.240000 324.820000 40.320000 ;
      RECT 236.620000 39.240000 279.820000 40.320000 ;
      RECT 191.620000 39.240000 234.820000 40.320000 ;
      RECT 146.620000 39.240000 189.820000 40.320000 ;
      RECT 101.620000 39.240000 144.820000 40.320000 ;
      RECT 56.620000 39.240000 99.820000 40.320000 ;
      RECT 11.620000 39.240000 54.820000 40.320000 ;
      RECT 4.860000 39.240000 9.655000 40.320000 ;
      RECT 0.000000 39.240000 2.260000 40.320000 ;
      RECT 0.000000 38.820000 548.960000 39.240000 ;
      RECT 0.000000 37.970000 550.160000 38.820000 ;
      RECT 0.000000 37.600000 548.960000 37.970000 ;
      RECT 544.900000 36.990000 548.960000 37.600000 ;
      RECT 544.900000 36.520000 550.160000 36.990000 ;
      RECT 508.620000 36.520000 542.300000 37.600000 ;
      RECT 463.620000 36.520000 506.820000 37.600000 ;
      RECT 418.620000 36.520000 461.820000 37.600000 ;
      RECT 373.620000 36.520000 416.820000 37.600000 ;
      RECT 328.620000 36.520000 371.820000 37.600000 ;
      RECT 283.620000 36.520000 326.820000 37.600000 ;
      RECT 238.620000 36.520000 281.820000 37.600000 ;
      RECT 193.620000 36.520000 236.820000 37.600000 ;
      RECT 148.620000 36.520000 191.820000 37.600000 ;
      RECT 103.620000 36.520000 146.820000 37.600000 ;
      RECT 58.620000 36.520000 101.820000 37.600000 ;
      RECT 13.620000 36.520000 56.820000 37.600000 ;
      RECT 7.860000 36.520000 11.820000 37.600000 ;
      RECT 0.000000 36.520000 5.260000 37.600000 ;
      RECT 0.000000 35.530000 550.160000 36.520000 ;
      RECT 0.000000 34.880000 548.960000 35.530000 ;
      RECT 547.900000 34.550000 548.960000 34.880000 ;
      RECT 547.900000 33.800000 550.160000 34.550000 ;
      RECT 506.620000 33.800000 545.300000 34.880000 ;
      RECT 461.620000 33.800000 504.820000 34.880000 ;
      RECT 416.620000 33.800000 459.820000 34.880000 ;
      RECT 371.620000 33.800000 414.820000 34.880000 ;
      RECT 326.620000 33.800000 369.820000 34.880000 ;
      RECT 281.620000 33.800000 324.820000 34.880000 ;
      RECT 236.620000 33.800000 279.820000 34.880000 ;
      RECT 191.620000 33.800000 234.820000 34.880000 ;
      RECT 146.620000 33.800000 189.820000 34.880000 ;
      RECT 101.620000 33.800000 144.820000 34.880000 ;
      RECT 56.620000 33.800000 99.820000 34.880000 ;
      RECT 11.620000 33.800000 54.820000 34.880000 ;
      RECT 4.860000 33.800000 9.655000 34.880000 ;
      RECT 0.000000 33.800000 2.260000 34.880000 ;
      RECT 0.000000 33.090000 550.160000 33.800000 ;
      RECT 0.000000 32.160000 548.960000 33.090000 ;
      RECT 544.900000 32.110000 548.960000 32.160000 ;
      RECT 544.900000 31.080000 550.160000 32.110000 ;
      RECT 508.620000 31.080000 542.300000 32.160000 ;
      RECT 463.620000 31.080000 506.820000 32.160000 ;
      RECT 418.620000 31.080000 461.820000 32.160000 ;
      RECT 373.620000 31.080000 416.820000 32.160000 ;
      RECT 328.620000 31.080000 371.820000 32.160000 ;
      RECT 283.620000 31.080000 326.820000 32.160000 ;
      RECT 238.620000 31.080000 281.820000 32.160000 ;
      RECT 193.620000 31.080000 236.820000 32.160000 ;
      RECT 148.620000 31.080000 191.820000 32.160000 ;
      RECT 103.620000 31.080000 146.820000 32.160000 ;
      RECT 58.620000 31.080000 101.820000 32.160000 ;
      RECT 13.620000 31.080000 56.820000 32.160000 ;
      RECT 7.860000 31.080000 11.820000 32.160000 ;
      RECT 0.000000 31.080000 5.260000 32.160000 ;
      RECT 0.000000 30.650000 550.160000 31.080000 ;
      RECT 0.000000 29.670000 548.960000 30.650000 ;
      RECT 0.000000 29.440000 550.160000 29.670000 ;
      RECT 547.900000 28.820000 550.160000 29.440000 ;
      RECT 547.900000 28.360000 548.960000 28.820000 ;
      RECT 506.620000 28.360000 545.300000 29.440000 ;
      RECT 461.620000 28.360000 504.820000 29.440000 ;
      RECT 416.620000 28.360000 459.820000 29.440000 ;
      RECT 371.620000 28.360000 414.820000 29.440000 ;
      RECT 326.620000 28.360000 369.820000 29.440000 ;
      RECT 281.620000 28.360000 324.820000 29.440000 ;
      RECT 236.620000 28.360000 279.820000 29.440000 ;
      RECT 191.620000 28.360000 234.820000 29.440000 ;
      RECT 146.620000 28.360000 189.820000 29.440000 ;
      RECT 101.620000 28.360000 144.820000 29.440000 ;
      RECT 56.620000 28.360000 99.820000 29.440000 ;
      RECT 11.620000 28.360000 54.820000 29.440000 ;
      RECT 4.860000 28.360000 9.655000 29.440000 ;
      RECT 0.000000 28.360000 2.260000 29.440000 ;
      RECT 0.000000 27.840000 548.960000 28.360000 ;
      RECT 0.000000 26.720000 550.160000 27.840000 ;
      RECT 544.900000 26.380000 550.160000 26.720000 ;
      RECT 544.900000 25.640000 548.960000 26.380000 ;
      RECT 508.620000 25.640000 542.300000 26.720000 ;
      RECT 463.620000 25.640000 506.820000 26.720000 ;
      RECT 418.620000 25.640000 461.820000 26.720000 ;
      RECT 373.620000 25.640000 416.820000 26.720000 ;
      RECT 328.620000 25.640000 371.820000 26.720000 ;
      RECT 283.620000 25.640000 326.820000 26.720000 ;
      RECT 238.620000 25.640000 281.820000 26.720000 ;
      RECT 193.620000 25.640000 236.820000 26.720000 ;
      RECT 148.620000 25.640000 191.820000 26.720000 ;
      RECT 103.620000 25.640000 146.820000 26.720000 ;
      RECT 58.620000 25.640000 101.820000 26.720000 ;
      RECT 13.620000 25.640000 56.820000 26.720000 ;
      RECT 7.860000 25.640000 11.820000 26.720000 ;
      RECT 0.000000 25.640000 5.260000 26.720000 ;
      RECT 0.000000 25.400000 548.960000 25.640000 ;
      RECT 0.000000 24.000000 550.160000 25.400000 ;
      RECT 547.900000 23.940000 550.160000 24.000000 ;
      RECT 547.900000 22.960000 548.960000 23.940000 ;
      RECT 547.900000 22.920000 550.160000 22.960000 ;
      RECT 506.620000 22.920000 545.300000 24.000000 ;
      RECT 461.620000 22.920000 504.820000 24.000000 ;
      RECT 416.620000 22.920000 459.820000 24.000000 ;
      RECT 371.620000 22.920000 414.820000 24.000000 ;
      RECT 326.620000 22.920000 369.820000 24.000000 ;
      RECT 281.620000 22.920000 324.820000 24.000000 ;
      RECT 236.620000 22.920000 279.820000 24.000000 ;
      RECT 191.620000 22.920000 234.820000 24.000000 ;
      RECT 146.620000 22.920000 189.820000 24.000000 ;
      RECT 101.620000 22.920000 144.820000 24.000000 ;
      RECT 56.620000 22.920000 99.820000 24.000000 ;
      RECT 11.620000 22.920000 54.820000 24.000000 ;
      RECT 4.860000 22.920000 9.655000 24.000000 ;
      RECT 0.000000 22.920000 2.260000 24.000000 ;
      RECT 0.000000 21.500000 550.160000 22.920000 ;
      RECT 0.000000 21.280000 548.960000 21.500000 ;
      RECT 544.900000 20.520000 548.960000 21.280000 ;
      RECT 544.900000 20.200000 550.160000 20.520000 ;
      RECT 508.620000 20.200000 542.300000 21.280000 ;
      RECT 463.620000 20.200000 506.820000 21.280000 ;
      RECT 418.620000 20.200000 461.820000 21.280000 ;
      RECT 373.620000 20.200000 416.820000 21.280000 ;
      RECT 328.620000 20.200000 371.820000 21.280000 ;
      RECT 283.620000 20.200000 326.820000 21.280000 ;
      RECT 238.620000 20.200000 281.820000 21.280000 ;
      RECT 193.620000 20.200000 236.820000 21.280000 ;
      RECT 148.620000 20.200000 191.820000 21.280000 ;
      RECT 103.620000 20.200000 146.820000 21.280000 ;
      RECT 58.620000 20.200000 101.820000 21.280000 ;
      RECT 13.620000 20.200000 56.820000 21.280000 ;
      RECT 7.860000 20.200000 11.820000 21.280000 ;
      RECT 0.000000 20.200000 5.260000 21.280000 ;
      RECT 0.000000 19.670000 550.160000 20.200000 ;
      RECT 0.000000 18.690000 548.960000 19.670000 ;
      RECT 0.000000 18.560000 550.160000 18.690000 ;
      RECT 547.900000 17.480000 550.160000 18.560000 ;
      RECT 506.620000 17.480000 545.300000 18.560000 ;
      RECT 461.620000 17.480000 504.820000 18.560000 ;
      RECT 416.620000 17.480000 459.820000 18.560000 ;
      RECT 371.620000 17.480000 414.820000 18.560000 ;
      RECT 326.620000 17.480000 369.820000 18.560000 ;
      RECT 281.620000 17.480000 324.820000 18.560000 ;
      RECT 236.620000 17.480000 279.820000 18.560000 ;
      RECT 191.620000 17.480000 234.820000 18.560000 ;
      RECT 146.620000 17.480000 189.820000 18.560000 ;
      RECT 101.620000 17.480000 144.820000 18.560000 ;
      RECT 56.620000 17.480000 99.820000 18.560000 ;
      RECT 11.620000 17.480000 54.820000 18.560000 ;
      RECT 4.860000 17.480000 9.655000 18.560000 ;
      RECT 0.000000 17.480000 2.260000 18.560000 ;
      RECT 0.000000 17.230000 550.160000 17.480000 ;
      RECT 0.000000 16.250000 548.960000 17.230000 ;
      RECT 0.000000 15.840000 550.160000 16.250000 ;
      RECT 544.900000 14.790000 550.160000 15.840000 ;
      RECT 544.900000 14.760000 548.960000 14.790000 ;
      RECT 508.620000 14.760000 542.300000 15.840000 ;
      RECT 463.620000 14.760000 506.820000 15.840000 ;
      RECT 418.620000 14.760000 461.820000 15.840000 ;
      RECT 373.620000 14.760000 416.820000 15.840000 ;
      RECT 328.620000 14.760000 371.820000 15.840000 ;
      RECT 283.620000 14.760000 326.820000 15.840000 ;
      RECT 238.620000 14.760000 281.820000 15.840000 ;
      RECT 193.620000 14.760000 236.820000 15.840000 ;
      RECT 148.620000 14.760000 191.820000 15.840000 ;
      RECT 103.620000 14.760000 146.820000 15.840000 ;
      RECT 58.620000 14.760000 101.820000 15.840000 ;
      RECT 13.620000 14.760000 56.820000 15.840000 ;
      RECT 7.860000 14.760000 11.820000 15.840000 ;
      RECT 0.000000 14.760000 5.260000 15.840000 ;
      RECT 0.000000 13.810000 548.960000 14.760000 ;
      RECT 0.000000 13.120000 550.160000 13.810000 ;
      RECT 547.900000 12.350000 550.160000 13.120000 ;
      RECT 547.900000 12.040000 548.960000 12.350000 ;
      RECT 506.620000 12.040000 545.300000 13.120000 ;
      RECT 461.620000 12.040000 504.820000 13.120000 ;
      RECT 416.620000 12.040000 459.820000 13.120000 ;
      RECT 371.620000 12.040000 414.820000 13.120000 ;
      RECT 326.620000 12.040000 369.820000 13.120000 ;
      RECT 281.620000 12.040000 324.820000 13.120000 ;
      RECT 236.620000 12.040000 279.820000 13.120000 ;
      RECT 191.620000 12.040000 234.820000 13.120000 ;
      RECT 146.620000 12.040000 189.820000 13.120000 ;
      RECT 101.620000 12.040000 144.820000 13.120000 ;
      RECT 56.620000 12.040000 99.820000 13.120000 ;
      RECT 11.620000 12.040000 54.820000 13.120000 ;
      RECT 4.860000 12.040000 9.655000 13.120000 ;
      RECT 0.000000 12.040000 2.260000 13.120000 ;
      RECT 0.000000 11.370000 548.960000 12.040000 ;
      RECT 0.000000 10.520000 550.160000 11.370000 ;
      RECT 0.000000 10.400000 548.960000 10.520000 ;
      RECT 544.900000 9.540000 548.960000 10.400000 ;
      RECT 544.900000 9.320000 550.160000 9.540000 ;
      RECT 508.620000 9.320000 542.300000 10.400000 ;
      RECT 463.620000 9.320000 506.820000 10.400000 ;
      RECT 418.620000 9.320000 461.820000 10.400000 ;
      RECT 373.620000 9.320000 416.820000 10.400000 ;
      RECT 328.620000 9.320000 371.820000 10.400000 ;
      RECT 283.620000 9.320000 326.820000 10.400000 ;
      RECT 238.620000 9.320000 281.820000 10.400000 ;
      RECT 193.620000 9.320000 236.820000 10.400000 ;
      RECT 148.620000 9.320000 191.820000 10.400000 ;
      RECT 103.620000 9.320000 146.820000 10.400000 ;
      RECT 58.620000 9.320000 101.820000 10.400000 ;
      RECT 13.620000 9.320000 56.820000 10.400000 ;
      RECT 7.860000 9.320000 11.820000 10.400000 ;
      RECT 0.000000 9.320000 5.260000 10.400000 ;
      RECT 0.000000 7.730000 550.160000 9.320000 ;
      RECT 0.000000 4.730000 550.160000 5.130000 ;
      RECT 0.000000 0.000000 550.160000 2.130000 ;
    LAYER met4 ;
      RECT 7.860000 546.460000 542.300000 549.780000 ;
      RECT 506.620000 543.460000 542.300000 546.460000 ;
      RECT 461.620000 543.460000 504.820000 546.460000 ;
      RECT 416.620000 543.460000 459.820000 546.460000 ;
      RECT 371.620000 543.460000 414.820000 546.460000 ;
      RECT 326.620000 543.460000 369.820000 546.460000 ;
      RECT 281.620000 543.460000 324.820000 546.460000 ;
      RECT 236.620000 543.460000 279.820000 546.460000 ;
      RECT 191.620000 543.460000 234.820000 546.460000 ;
      RECT 146.620000 543.460000 189.820000 546.460000 ;
      RECT 101.620000 543.460000 144.820000 546.460000 ;
      RECT 56.620000 543.460000 99.820000 546.460000 ;
      RECT 11.620000 543.460000 54.820000 546.460000 ;
      RECT 7.860000 535.360000 9.820000 546.460000 ;
      RECT 7.860000 534.280000 9.655000 535.360000 ;
      RECT 7.860000 529.920000 9.820000 534.280000 ;
      RECT 7.860000 528.840000 9.655000 529.920000 ;
      RECT 7.860000 524.480000 9.820000 528.840000 ;
      RECT 7.860000 523.400000 9.655000 524.480000 ;
      RECT 7.860000 519.040000 9.820000 523.400000 ;
      RECT 7.860000 517.960000 9.655000 519.040000 ;
      RECT 7.860000 513.600000 9.820000 517.960000 ;
      RECT 7.860000 512.520000 9.655000 513.600000 ;
      RECT 7.860000 508.160000 9.820000 512.520000 ;
      RECT 7.860000 507.080000 9.655000 508.160000 ;
      RECT 7.860000 502.720000 9.820000 507.080000 ;
      RECT 7.860000 501.640000 9.655000 502.720000 ;
      RECT 7.860000 497.280000 9.820000 501.640000 ;
      RECT 7.860000 496.200000 9.655000 497.280000 ;
      RECT 7.860000 491.840000 9.820000 496.200000 ;
      RECT 7.860000 490.760000 9.655000 491.840000 ;
      RECT 7.860000 486.400000 9.820000 490.760000 ;
      RECT 7.860000 485.320000 9.655000 486.400000 ;
      RECT 7.860000 480.960000 9.820000 485.320000 ;
      RECT 7.860000 479.880000 9.655000 480.960000 ;
      RECT 7.860000 475.520000 9.820000 479.880000 ;
      RECT 7.860000 474.440000 9.655000 475.520000 ;
      RECT 7.860000 470.080000 9.820000 474.440000 ;
      RECT 7.860000 469.000000 9.655000 470.080000 ;
      RECT 7.860000 464.640000 9.820000 469.000000 ;
      RECT 7.860000 463.560000 9.655000 464.640000 ;
      RECT 7.860000 459.200000 9.820000 463.560000 ;
      RECT 7.860000 458.120000 9.655000 459.200000 ;
      RECT 7.860000 453.760000 9.820000 458.120000 ;
      RECT 7.860000 452.680000 9.655000 453.760000 ;
      RECT 7.860000 448.320000 9.820000 452.680000 ;
      RECT 7.860000 447.240000 9.655000 448.320000 ;
      RECT 7.860000 442.880000 9.820000 447.240000 ;
      RECT 7.860000 441.800000 9.655000 442.880000 ;
      RECT 7.860000 437.440000 9.820000 441.800000 ;
      RECT 7.860000 436.360000 9.655000 437.440000 ;
      RECT 7.860000 432.000000 9.820000 436.360000 ;
      RECT 7.860000 430.920000 9.655000 432.000000 ;
      RECT 7.860000 426.560000 9.820000 430.920000 ;
      RECT 7.860000 425.480000 9.655000 426.560000 ;
      RECT 7.860000 421.120000 9.820000 425.480000 ;
      RECT 7.860000 420.040000 9.655000 421.120000 ;
      RECT 7.860000 415.680000 9.820000 420.040000 ;
      RECT 7.860000 414.600000 9.655000 415.680000 ;
      RECT 7.860000 410.240000 9.820000 414.600000 ;
      RECT 7.860000 409.160000 9.655000 410.240000 ;
      RECT 7.860000 404.800000 9.820000 409.160000 ;
      RECT 7.860000 403.720000 9.655000 404.800000 ;
      RECT 7.860000 399.360000 9.820000 403.720000 ;
      RECT 7.860000 398.280000 9.655000 399.360000 ;
      RECT 7.860000 393.920000 9.820000 398.280000 ;
      RECT 7.860000 392.840000 9.655000 393.920000 ;
      RECT 7.860000 388.480000 9.820000 392.840000 ;
      RECT 7.860000 387.400000 9.655000 388.480000 ;
      RECT 7.860000 383.040000 9.820000 387.400000 ;
      RECT 7.860000 381.960000 9.655000 383.040000 ;
      RECT 7.860000 377.600000 9.820000 381.960000 ;
      RECT 7.860000 376.520000 9.655000 377.600000 ;
      RECT 7.860000 372.160000 9.820000 376.520000 ;
      RECT 7.860000 371.080000 9.655000 372.160000 ;
      RECT 7.860000 366.720000 9.820000 371.080000 ;
      RECT 7.860000 365.640000 9.655000 366.720000 ;
      RECT 7.860000 361.280000 9.820000 365.640000 ;
      RECT 7.860000 360.200000 9.655000 361.280000 ;
      RECT 7.860000 355.840000 9.820000 360.200000 ;
      RECT 7.860000 354.760000 9.655000 355.840000 ;
      RECT 7.860000 350.400000 9.820000 354.760000 ;
      RECT 7.860000 349.320000 9.655000 350.400000 ;
      RECT 7.860000 344.960000 9.820000 349.320000 ;
      RECT 7.860000 343.880000 9.655000 344.960000 ;
      RECT 7.860000 339.520000 9.820000 343.880000 ;
      RECT 7.860000 338.440000 9.655000 339.520000 ;
      RECT 7.860000 334.080000 9.820000 338.440000 ;
      RECT 7.860000 333.000000 9.655000 334.080000 ;
      RECT 7.860000 328.640000 9.820000 333.000000 ;
      RECT 7.860000 327.560000 9.655000 328.640000 ;
      RECT 7.860000 323.200000 9.820000 327.560000 ;
      RECT 7.860000 322.120000 9.655000 323.200000 ;
      RECT 7.860000 317.760000 9.820000 322.120000 ;
      RECT 7.860000 316.680000 9.655000 317.760000 ;
      RECT 7.860000 312.320000 9.820000 316.680000 ;
      RECT 7.860000 311.240000 9.655000 312.320000 ;
      RECT 7.860000 306.880000 9.820000 311.240000 ;
      RECT 7.860000 305.800000 9.655000 306.880000 ;
      RECT 7.860000 301.440000 9.820000 305.800000 ;
      RECT 7.860000 300.360000 9.655000 301.440000 ;
      RECT 7.860000 296.000000 9.820000 300.360000 ;
      RECT 7.860000 294.920000 9.655000 296.000000 ;
      RECT 7.860000 290.560000 9.820000 294.920000 ;
      RECT 7.860000 289.480000 9.655000 290.560000 ;
      RECT 7.860000 285.120000 9.820000 289.480000 ;
      RECT 7.860000 284.040000 9.655000 285.120000 ;
      RECT 7.860000 279.680000 9.820000 284.040000 ;
      RECT 7.860000 278.600000 9.655000 279.680000 ;
      RECT 7.860000 274.240000 9.820000 278.600000 ;
      RECT 7.860000 273.160000 9.655000 274.240000 ;
      RECT 7.860000 268.800000 9.820000 273.160000 ;
      RECT 7.860000 267.720000 9.655000 268.800000 ;
      RECT 7.860000 263.360000 9.820000 267.720000 ;
      RECT 7.860000 262.280000 9.655000 263.360000 ;
      RECT 7.860000 257.920000 9.820000 262.280000 ;
      RECT 7.860000 256.840000 9.655000 257.920000 ;
      RECT 7.860000 252.480000 9.820000 256.840000 ;
      RECT 7.860000 251.400000 9.655000 252.480000 ;
      RECT 7.860000 247.040000 9.820000 251.400000 ;
      RECT 7.860000 245.960000 9.655000 247.040000 ;
      RECT 7.860000 241.600000 9.820000 245.960000 ;
      RECT 7.860000 240.520000 9.655000 241.600000 ;
      RECT 7.860000 236.160000 9.820000 240.520000 ;
      RECT 7.860000 235.080000 9.655000 236.160000 ;
      RECT 7.860000 230.720000 9.820000 235.080000 ;
      RECT 7.860000 229.640000 9.655000 230.720000 ;
      RECT 7.860000 225.280000 9.820000 229.640000 ;
      RECT 7.860000 224.200000 9.655000 225.280000 ;
      RECT 7.860000 219.840000 9.820000 224.200000 ;
      RECT 7.860000 218.760000 9.655000 219.840000 ;
      RECT 7.860000 214.400000 9.820000 218.760000 ;
      RECT 7.860000 213.320000 9.655000 214.400000 ;
      RECT 7.860000 208.960000 9.820000 213.320000 ;
      RECT 7.860000 207.880000 9.655000 208.960000 ;
      RECT 7.860000 203.520000 9.820000 207.880000 ;
      RECT 7.860000 202.440000 9.655000 203.520000 ;
      RECT 7.860000 198.080000 9.820000 202.440000 ;
      RECT 7.860000 197.000000 9.655000 198.080000 ;
      RECT 7.860000 192.640000 9.820000 197.000000 ;
      RECT 7.860000 191.560000 9.655000 192.640000 ;
      RECT 7.860000 187.200000 9.820000 191.560000 ;
      RECT 7.860000 186.120000 9.655000 187.200000 ;
      RECT 7.860000 181.760000 9.820000 186.120000 ;
      RECT 7.860000 180.680000 9.655000 181.760000 ;
      RECT 7.860000 176.320000 9.820000 180.680000 ;
      RECT 7.860000 175.240000 9.655000 176.320000 ;
      RECT 7.860000 170.880000 9.820000 175.240000 ;
      RECT 7.860000 169.800000 9.655000 170.880000 ;
      RECT 7.860000 165.440000 9.820000 169.800000 ;
      RECT 7.860000 164.360000 9.655000 165.440000 ;
      RECT 7.860000 160.000000 9.820000 164.360000 ;
      RECT 7.860000 158.920000 9.655000 160.000000 ;
      RECT 7.860000 154.560000 9.820000 158.920000 ;
      RECT 7.860000 153.480000 9.655000 154.560000 ;
      RECT 7.860000 149.120000 9.820000 153.480000 ;
      RECT 7.860000 148.040000 9.655000 149.120000 ;
      RECT 7.860000 143.680000 9.820000 148.040000 ;
      RECT 7.860000 142.600000 9.655000 143.680000 ;
      RECT 7.860000 138.240000 9.820000 142.600000 ;
      RECT 7.860000 137.160000 9.655000 138.240000 ;
      RECT 7.860000 132.800000 9.820000 137.160000 ;
      RECT 7.860000 131.720000 9.655000 132.800000 ;
      RECT 7.860000 127.360000 9.820000 131.720000 ;
      RECT 7.860000 126.280000 9.655000 127.360000 ;
      RECT 7.860000 121.920000 9.820000 126.280000 ;
      RECT 7.860000 120.840000 9.655000 121.920000 ;
      RECT 7.860000 116.480000 9.820000 120.840000 ;
      RECT 7.860000 115.400000 9.655000 116.480000 ;
      RECT 7.860000 111.040000 9.820000 115.400000 ;
      RECT 7.860000 109.960000 9.655000 111.040000 ;
      RECT 7.860000 105.600000 9.820000 109.960000 ;
      RECT 7.860000 104.520000 9.655000 105.600000 ;
      RECT 7.860000 100.160000 9.820000 104.520000 ;
      RECT 7.860000 99.080000 9.655000 100.160000 ;
      RECT 7.860000 94.720000 9.820000 99.080000 ;
      RECT 7.860000 93.640000 9.655000 94.720000 ;
      RECT 7.860000 89.280000 9.820000 93.640000 ;
      RECT 7.860000 88.200000 9.655000 89.280000 ;
      RECT 7.860000 83.840000 9.820000 88.200000 ;
      RECT 7.860000 82.760000 9.655000 83.840000 ;
      RECT 7.860000 78.400000 9.820000 82.760000 ;
      RECT 7.860000 77.320000 9.655000 78.400000 ;
      RECT 7.860000 72.960000 9.820000 77.320000 ;
      RECT 7.860000 71.880000 9.655000 72.960000 ;
      RECT 7.860000 67.520000 9.820000 71.880000 ;
      RECT 7.860000 66.440000 9.655000 67.520000 ;
      RECT 7.860000 62.080000 9.820000 66.440000 ;
      RECT 7.860000 61.000000 9.655000 62.080000 ;
      RECT 7.860000 56.640000 9.820000 61.000000 ;
      RECT 7.860000 55.560000 9.655000 56.640000 ;
      RECT 7.860000 51.200000 9.820000 55.560000 ;
      RECT 7.860000 50.120000 9.655000 51.200000 ;
      RECT 7.860000 45.760000 9.820000 50.120000 ;
      RECT 7.860000 44.680000 9.655000 45.760000 ;
      RECT 7.860000 40.320000 9.820000 44.680000 ;
      RECT 7.860000 39.240000 9.655000 40.320000 ;
      RECT 7.860000 34.880000 9.820000 39.240000 ;
      RECT 7.860000 33.800000 9.655000 34.880000 ;
      RECT 7.860000 29.440000 9.820000 33.800000 ;
      RECT 7.860000 28.360000 9.655000 29.440000 ;
      RECT 7.860000 24.000000 9.820000 28.360000 ;
      RECT 7.860000 22.920000 9.655000 24.000000 ;
      RECT 7.860000 18.560000 9.820000 22.920000 ;
      RECT 7.860000 17.480000 9.655000 18.560000 ;
      RECT 7.860000 13.120000 9.820000 17.480000 ;
      RECT 7.860000 12.040000 9.655000 13.120000 ;
      RECT 508.620000 5.130000 542.300000 543.460000 ;
      RECT 506.620000 5.130000 506.820000 543.460000 ;
      RECT 463.620000 5.130000 504.820000 543.460000 ;
      RECT 461.620000 5.130000 461.820000 543.460000 ;
      RECT 418.620000 5.130000 459.820000 543.460000 ;
      RECT 416.620000 5.130000 416.820000 543.460000 ;
      RECT 373.620000 5.130000 414.820000 543.460000 ;
      RECT 371.620000 5.130000 371.820000 543.460000 ;
      RECT 328.620000 5.130000 369.820000 543.460000 ;
      RECT 326.620000 5.130000 326.820000 543.460000 ;
      RECT 283.620000 5.130000 324.820000 543.460000 ;
      RECT 281.620000 5.130000 281.820000 543.460000 ;
      RECT 238.620000 5.130000 279.820000 543.460000 ;
      RECT 236.620000 5.130000 236.820000 543.460000 ;
      RECT 193.620000 5.130000 234.820000 543.460000 ;
      RECT 191.620000 5.130000 191.820000 543.460000 ;
      RECT 148.620000 5.130000 189.820000 543.460000 ;
      RECT 146.620000 5.130000 146.820000 543.460000 ;
      RECT 103.620000 5.130000 144.820000 543.460000 ;
      RECT 101.620000 5.130000 101.820000 543.460000 ;
      RECT 58.620000 5.130000 99.820000 543.460000 ;
      RECT 56.620000 5.130000 56.820000 543.460000 ;
      RECT 13.620000 5.130000 54.820000 543.460000 ;
      RECT 11.620000 5.130000 11.820000 543.460000 ;
      RECT 506.620000 2.130000 542.300000 5.130000 ;
      RECT 461.620000 2.130000 504.820000 5.130000 ;
      RECT 416.620000 2.130000 459.820000 5.130000 ;
      RECT 371.620000 2.130000 414.820000 5.130000 ;
      RECT 326.620000 2.130000 369.820000 5.130000 ;
      RECT 281.620000 2.130000 324.820000 5.130000 ;
      RECT 236.620000 2.130000 279.820000 5.130000 ;
      RECT 191.620000 2.130000 234.820000 5.130000 ;
      RECT 146.620000 2.130000 189.820000 5.130000 ;
      RECT 101.620000 2.130000 144.820000 5.130000 ;
      RECT 56.620000 2.130000 99.820000 5.130000 ;
      RECT 11.620000 2.130000 54.820000 5.130000 ;
      RECT 7.860000 2.130000 9.820000 12.040000 ;
      RECT 547.900000 0.000000 550.160000 549.780000 ;
      RECT 544.900000 0.000000 545.300000 549.780000 ;
      RECT 7.860000 0.000000 542.300000 2.130000 ;
      RECT 4.860000 0.000000 5.260000 549.780000 ;
      RECT 0.000000 0.000000 2.260000 549.780000 ;
  END
END ibex_core

END LIBRARY
