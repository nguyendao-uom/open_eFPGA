##
## LEF for PtnCells ;
## created by Innovus v19.11-s128_1 on Thu Dec 23 11:05:55 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO ibex_top
  CLASS BLOCK ;
  SIZE 550.160000 BY 599.760000 ;
  FOREIGN ibex_top 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.4456 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.984 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.304 LAYER met3  ;
    ANTENNAMAXAREACAR 1.8071 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 7.68359 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.0396701 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 10.160000 0.000000 10.540000 0.900000 ;
    END
  END clk_i
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1851 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.6554 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.84 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 7.8795 LAYER met3  ;
    ANTENNAMAXAREACAR 28.2255 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 137.482 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.678855 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 40.2759 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 217.152 LAYER met4  ;
    ANTENNAGATEAREA 13.2495 LAYER met4  ;
    ANTENNAMAXAREACAR 31.2653 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 153.871 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.678855 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 11.080000 0.000000 11.460000 0.900000 ;
    END
  END rst_ni
  PIN test_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9438 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.611 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 20.1444 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 91.6786 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 12.460000 0.000000 12.840000 0.900000 ;
    END
  END test_en_i
  PIN ram_cfg_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.840000 0.000000 14.220000 0.900000 ;
    END
  END ram_cfg_i
  PIN hart_id_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.3336 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.3258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 18.5111 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 96.0323 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 15.220000 0.000000 15.600000 0.900000 ;
    END
  END hart_id_i[31]
  PIN hart_id_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1387 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.2965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.0782 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.632 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 66.322 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 352.032 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 16.140000 0.000000 16.520000 0.900000 ;
    END
  END hart_id_i[30]
  PIN hart_id_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.1707 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.6925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.6608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.328 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 45.5154 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 235.398 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 17.520000 0.000000 17.900000 0.900000 ;
    END
  END hart_id_i[29]
  PIN hart_id_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.5237 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.4575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.9388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.144 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 51.7501 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 273.083 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 18.900000 0.000000 19.280000 0.900000 ;
    END
  END hart_id_i[28]
  PIN hart_id_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.1993 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.7175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.7388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.744 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 65.9226 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 342.057 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 20.280000 0.000000 20.660000 0.900000 ;
    END
  END hart_id_i[27]
  PIN hart_id_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6121 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.0138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 96.544 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 111.234 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 591.636 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 21.660000 0.000000 22.040000 0.900000 ;
    END
  END hart_id_i[26]
  PIN hart_id_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6121 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.286 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.1248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 81.136 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 77.0034 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 409.968 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 22.580000 0.000000 22.960000 0.900000 ;
    END
  END hart_id_i[25]
  PIN hart_id_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4413 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.8418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 84.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 110.427 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 586.941 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 23.960000 0.000000 24.340000 0.900000 ;
    END
  END hart_id_i[24]
  PIN hart_id_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.7626 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.587 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 40.6952 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 199.606 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 25.340000 0.000000 25.720000 0.900000 ;
    END
  END hart_id_i[23]
  PIN hart_id_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9097 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.1515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.1736 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 55.2956 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 290.061 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 26.720000 0.000000 27.100000 0.900000 ;
    END
  END hart_id_i[22]
  PIN hart_id_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.9593 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 89.2815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.6996 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.672 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 69.138 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 362.448 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 27.640000 0.000000 28.020000 0.900000 ;
    END
  END hart_id_i[21]
  PIN hart_id_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7977 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.7095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.4206 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.984 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 19.4117 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 103.739 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 29.020000 0.000000 29.400000 0.900000 ;
    END
  END hart_id_i[20]
  PIN hart_id_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.3861 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.4155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.0236 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.4 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 66.6467 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 350.655 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 30.400000 0.000000 30.780000 0.900000 ;
    END
  END hart_id_i[19]
  PIN hart_id_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7517 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.3615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.3116 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.936 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 53.2002 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 279.77 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 31.780000 0.000000 32.160000 0.900000 ;
    END
  END hart_id_i[18]
  PIN hart_id_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8763 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.1025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 32.7604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 176.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 17.0103 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 90.9899 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 33.160000 0.000000 33.540000 0.900000 ;
    END
  END hart_id_i[17]
  PIN hart_id_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.3755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.3952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.656 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 26.0319 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 140.711 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 34.080000 0.000000 34.460000 0.900000 ;
    END
  END hart_id_i[16]
  PIN hart_id_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.1697 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.5695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.1846 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 52.1541 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 274.848 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 35.460000 0.000000 35.840000 0.900000 ;
    END
  END hart_id_i[15]
  PIN hart_id_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0483 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.9625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.4184 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.976 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 56.7576 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 304.493 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 36.840000 0.000000 37.220000 0.900000 ;
    END
  END hart_id_i[14]
  PIN hart_id_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7055 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.2485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.3542 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.104 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 63.7143 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 340.271 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 38.220000 0.000000 38.600000 0.900000 ;
    END
  END hart_id_i[13]
  PIN hart_id_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9537 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.2138 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 52.3616 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 285.135 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 39.140000 0.000000 39.520000 0.900000 ;
    END
  END hart_id_i[12]
  PIN hart_id_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0143 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 32.0956 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 172.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 9.12727 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 50.1535 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 40.520000 0.000000 40.900000 0.900000 ;
    END
  END hart_id_i[11]
  PIN hart_id_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6307 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.5205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.2124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 72.9665 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 388.008 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 41.900000 0.000000 42.280000 0.900000 ;
    END
  END hart_id_i[10]
  PIN hart_id_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.394 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.13838 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.9859 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 43.280000 0.000000 43.660000 0.900000 ;
    END
  END hart_id_i[9]
  PIN hart_id_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.8352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 148.897 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.9728 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.992 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 25.8982 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 136.149 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 44.660000 0.000000 45.040000 0.900000 ;
    END
  END hart_id_i[8]
  PIN hart_id_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.9758 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 128.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 43.3572 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 229.834 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 45.580000 0.000000 45.960000 0.900000 ;
    END
  END hart_id_i[7]
  PIN hart_id_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5057 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.6788 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 15.8089 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 83.6404 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 46.960000 0.000000 47.340000 0.900000 ;
    END
  END hart_id_i[6]
  PIN hart_id_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5949 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.9988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 150.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 23.6218 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 125.2 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 48.340000 0.000000 48.720000 0.900000 ;
    END
  END hart_id_i[5]
  PIN hart_id_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0395 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.9185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.77 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.792 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 40.4865 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 218.784 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 49.720000 0.000000 50.100000 0.900000 ;
    END
  END hart_id_i[4]
  PIN hart_id_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.9275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.3188 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 17.1354 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 90.4606 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 50.640000 0.000000 51.020000 0.900000 ;
    END
  END hart_id_i[3]
  PIN hart_id_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.6349 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.0135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.1764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 138.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.8846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.992 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 24.5002 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 131.37 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 52.020000 0.000000 52.400000 0.900000 ;
    END
  END hart_id_i[2]
  PIN hart_id_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0143 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.8724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 171.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 11.2473 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 61.8505 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 53.400000 0.000000 53.780000 0.900000 ;
    END
  END hart_id_i[1]
  PIN hart_id_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5539 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.3725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.3816 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.976 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 65.6877 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 344.562 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 54.780000 0.000000 55.160000 0.900000 ;
    END
  END hart_id_i[0]
  PIN boot_addr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5419 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.9626 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.408 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 82.1968 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 417.034 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 56.160000 0.000000 56.540000 0.900000 ;
    END
  END boot_addr_i[31]
  PIN boot_addr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0787 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.1248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 81.136 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 108.065 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 553.329 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 57.080000 0.000000 57.460000 0.900000 ;
    END
  END boot_addr_i[30]
  PIN boot_addr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4413 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.4778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 72.352 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 105.186 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 533.76 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 58.460000 0.000000 58.840000 0.900000 ;
    END
  END boot_addr_i[29]
  PIN boot_addr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2609 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.1435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.471 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.3604 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 78 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 103.206 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 534.845 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.67778 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 59.840000 0.000000 60.220000 0.900000 ;
    END
  END boot_addr_i[28]
  PIN boot_addr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4207 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.229 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.1948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.176 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 61.1885 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 301.585 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 61.220000 0.000000 61.600000 0.900000 ;
    END
  END boot_addr_i[27]
  PIN boot_addr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4413 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.5148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 83.216 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 83.5357 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 424.202 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 62.140000 0.000000 62.520000 0.900000 ;
    END
  END boot_addr_i[26]
  PIN boot_addr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.373 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 41.754 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 190.135 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 63.520000 0.000000 63.900000 0.900000 ;
    END
  END boot_addr_i[25]
  PIN boot_addr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4847 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.3058 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 76.768 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 80.1694 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 406.776 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 64.900000 0.000000 65.280000 0.900000 ;
    END
  END boot_addr_i[24]
  PIN boot_addr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3425 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.3778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 45.152 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 56.6321 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 279.514 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 66.280000 0.000000 66.660000 0.900000 ;
    END
  END boot_addr_i[23]
  PIN boot_addr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0143 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.2818 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 76.64 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 77.6893 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 393.613 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 67.660000 0.000000 68.040000 0.900000 ;
    END
  END boot_addr_i[22]
  PIN boot_addr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8339 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.0085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.056 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.2558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.168 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 48.7012 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 238.649 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 68.580000 0.000000 68.960000 0.900000 ;
    END
  END boot_addr_i[21]
  PIN boot_addr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5949 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.1838 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 54.784 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 82.9401 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 421.153 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 69.960000 0.000000 70.340000 0.900000 ;
    END
  END boot_addr_i[20]
  PIN boot_addr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2385 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.0315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.953 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.2188 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.304 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 48.8413 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 240.385 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 71.340000 0.000000 71.720000 0.900000 ;
    END
  END boot_addr_i[19]
  PIN boot_addr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.3865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.7808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 57.968 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 63.5742 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 318.407 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 72.720000 0.000000 73.100000 0.900000 ;
    END
  END boot_addr_i[18]
  PIN boot_addr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.5215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.4148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 56.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 75.8139 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 382.395 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 74.100000 0.000000 74.480000 0.900000 ;
    END
  END boot_addr_i[17]
  PIN boot_addr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.801 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.1598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.656 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 82.4623 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 416.815 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 75.020000 0.000000 75.400000 0.900000 ;
    END
  END boot_addr_i[16]
  PIN boot_addr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3559 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.619 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.8808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 85.168 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 90.0095 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 459.496 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 76.400000 0.000000 76.780000 0.900000 ;
    END
  END boot_addr_i[15]
  PIN boot_addr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7289 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.4835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.8548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 63.696 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 97.5786 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 499.52 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 77.780000 0.000000 78.160000 0.900000 ;
    END
  END boot_addr_i[14]
  PIN boot_addr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2537 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.9895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.0838 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.584 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 80.8321 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 401.74 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 79.160000 0.000000 79.540000 0.900000 ;
    END
  END boot_addr_i[13]
  PIN boot_addr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.1086 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 81.52 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 108.465 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 550.331 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 80.080000 0.000000 80.460000 0.900000 ;
    END
  END boot_addr_i[12]
  PIN boot_addr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7619 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.963 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.8418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 68.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 92.5909 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 468.942 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 81.460000 0.000000 81.840000 0.900000 ;
    END
  END boot_addr_i[11]
  PIN boot_addr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6861 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.677 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.3156 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 98.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 115.727 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 591.103 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.85635 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 82.840000 0.000000 83.220000 0.900000 ;
    END
  END boot_addr_i[10]
  PIN boot_addr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.056 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.1098 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 65.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 129.073 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 649.579 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.884127 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 84.220000 0.000000 84.600000 0.900000 ;
    END
  END boot_addr_i[9]
  PIN boot_addr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.736 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.392 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.5868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 83.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 129.171 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 654.885 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.20159 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 85.600000 0.000000 85.980000 0.900000 ;
    END
  END boot_addr_i[8]
  PIN boot_addr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.520000 0.000000 86.900000 0.900000 ;
    END
  END boot_addr_i[7]
  PIN boot_addr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.900000 0.000000 88.280000 0.900000 ;
    END
  END boot_addr_i[6]
  PIN boot_addr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.280000 0.000000 89.660000 0.900000 ;
    END
  END boot_addr_i[5]
  PIN boot_addr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.660000 0.000000 91.040000 0.900000 ;
    END
  END boot_addr_i[4]
  PIN boot_addr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.580000 0.000000 91.960000 0.900000 ;
    END
  END boot_addr_i[3]
  PIN boot_addr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.960000 0.000000 93.340000 0.900000 ;
    END
  END boot_addr_i[2]
  PIN boot_addr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.340000 0.000000 94.720000 0.900000 ;
    END
  END boot_addr_i[1]
  PIN boot_addr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.720000 0.000000 96.100000 0.900000 ;
    END
  END boot_addr_i[0]
  PIN instr_req_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1773 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.04072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.664 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 97.100000 0.000000 97.480000 0.900000 ;
    END
  END instr_req_o
  PIN instr_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5016 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.39 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 22.6004 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 108.29 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 98.020000 0.000000 98.400000 0.900000 ;
    END
  END instr_gnt_i
  PIN instr_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0696 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.122 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 13.2576 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.7919 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 99.400000 0.000000 99.780000 0.900000 ;
    END
  END instr_rvalid_i
  PIN instr_addr_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2966 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.375 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 100.780000 0.000000 101.160000 0.900000 ;
    END
  END instr_addr_o[31]
  PIN instr_addr_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7798 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.673 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 102.160000 0.000000 102.540000 0.900000 ;
    END
  END instr_addr_o[30]
  PIN instr_addr_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9842 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.695 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 103.080000 0.000000 103.460000 0.900000 ;
    END
  END instr_addr_o[29]
  PIN instr_addr_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.001 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.779 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 104.460000 0.000000 104.840000 0.900000 ;
    END
  END instr_addr_o[28]
  PIN instr_addr_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6982 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.265 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 105.840000 0.000000 106.220000 0.900000 ;
    END
  END instr_addr_o[27]
  PIN instr_addr_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6034 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.791 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 107.220000 0.000000 107.600000 0.900000 ;
    END
  END instr_addr_o[26]
  PIN instr_addr_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5558 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.553 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 108.600000 0.000000 108.980000 0.900000 ;
    END
  END instr_addr_o[25]
  PIN instr_addr_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0486 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.017 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 109.520000 0.000000 109.900000 0.900000 ;
    END
  END instr_addr_o[24]
  PIN instr_addr_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6244 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.896 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 110.900000 0.000000 111.280000 0.900000 ;
    END
  END instr_addr_o[23]
  PIN instr_addr_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.106 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 112.280000 0.000000 112.660000 0.900000 ;
    END
  END instr_addr_o[22]
  PIN instr_addr_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6034 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.791 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 113.660000 0.000000 114.040000 0.900000 ;
    END
  END instr_addr_o[21]
  PIN instr_addr_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4646 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.215 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 114.580000 0.000000 114.960000 0.900000 ;
    END
  END instr_addr_o[20]
  PIN instr_addr_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.599 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 115.960000 0.000000 116.340000 0.900000 ;
    END
  END instr_addr_o[19]
  PIN instr_addr_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 117.340000 0.000000 117.720000 0.900000 ;
    END
  END instr_addr_o[18]
  PIN instr_addr_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.529 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.537 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 118.720000 0.000000 119.100000 0.900000 ;
    END
  END instr_addr_o[17]
  PIN instr_addr_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8006 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.895 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 120.100000 0.000000 120.480000 0.900000 ;
    END
  END instr_addr_o[16]
  PIN instr_addr_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.435 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 121.020000 0.000000 121.400000 0.900000 ;
    END
  END instr_addr_o[15]
  PIN instr_addr_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4342 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.063 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 122.400000 0.000000 122.780000 0.900000 ;
    END
  END instr_addr_o[14]
  PIN instr_addr_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7092 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.428 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 123.780000 0.000000 124.160000 0.900000 ;
    END
  END instr_addr_o[13]
  PIN instr_addr_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.563 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.707 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 125.160000 0.000000 125.540000 0.900000 ;
    END
  END instr_addr_o[12]
  PIN instr_addr_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4366 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.075 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 126.080000 0.000000 126.460000 0.900000 ;
    END
  END instr_addr_o[11]
  PIN instr_addr_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.435 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 127.460000 0.000000 127.840000 0.900000 ;
    END
  END instr_addr_o[10]
  PIN instr_addr_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.729 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 128.840000 0.000000 129.220000 0.900000 ;
    END
  END instr_addr_o[9]
  PIN instr_addr_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.651 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.029 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 130.220000 0.000000 130.600000 0.900000 ;
    END
  END instr_addr_o[8]
  PIN instr_addr_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7362 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 131.600000 0.000000 131.980000 0.900000 ;
    END
  END instr_addr_o[7]
  PIN instr_addr_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.389 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.837 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 132.520000 0.000000 132.900000 0.900000 ;
    END
  END instr_addr_o[6]
  PIN instr_addr_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4818 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.301 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 133.900000 0.000000 134.280000 0.900000 ;
    END
  END instr_addr_o[5]
  PIN instr_addr_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8274 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.911 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 135.280000 0.000000 135.660000 0.900000 ;
    END
  END instr_addr_o[4]
  PIN instr_addr_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6121 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.2248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.336 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 136.660000 0.000000 137.040000 0.900000 ;
    END
  END instr_addr_o[3]
  PIN instr_addr_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.599 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 138.040000 0.000000 138.420000 0.900000 ;
    END
  END instr_addr_o[2]
  PIN instr_addr_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.889 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.219 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 138.960000 0.000000 139.340000 0.900000 ;
    END
  END instr_addr_o[1]
  PIN instr_addr_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.563 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.707 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 140.340000 0.000000 140.720000 0.900000 ;
    END
  END instr_addr_o[0]
  PIN instr_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4847 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.446 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.0488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 54.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6255 LAYER met4  ;
    ANTENNAMAXAREACAR 46.7655 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 230.888 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.756277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 141.720000 0.000000 142.100000 0.900000 ;
    END
  END instr_rdata_i[31]
  PIN instr_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.9758 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.319 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6255 LAYER met2  ;
    ANTENNAMAXAREACAR 24.0515 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 108.34 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 143.100000 0.000000 143.480000 0.900000 ;
    END
  END instr_rdata_i[30]
  PIN instr_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.1818 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 49.44 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6255 LAYER met4  ;
    ANTENNAMAXAREACAR 28.4068 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 136.623 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.535834 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 144.020000 0.000000 144.400000 0.900000 ;
    END
  END instr_rdata_i[29]
  PIN instr_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.1994 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.535 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6255 LAYER met2  ;
    ANTENNAMAXAREACAR 30.8553 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 142.195 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 145.400000 0.000000 145.780000 0.900000 ;
    END
  END instr_rdata_i[28]
  PIN instr_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9669 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.2215 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4995 LAYER met2  ;
    ANTENNAMAXAREACAR 20.9573 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 92.5372 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.488017 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.6378 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.872 LAYER met3  ;
    ANTENNAGATEAREA 0.6255 LAYER met3  ;
    ANTENNAMAXAREACAR 36.3654 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 175.466 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 146.780000 0.000000 147.160000 0.900000 ;
    END
  END instr_rdata_i[27]
  PIN instr_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.383 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6255 LAYER met2  ;
    ANTENNAMAXAREACAR 17.8201 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.1836 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 148.160000 0.000000 148.540000 0.900000 ;
    END
  END instr_rdata_i[26]
  PIN instr_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7697 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.2255 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 LAYER met2  ;
    ANTENNAMAXAREACAR 37.2573 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 173.295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.692328 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met3  ;
    ANTENNAGATEAREA 0.6255 LAYER met3  ;
    ANTENNAMAXAREACAR 39.4328 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 185.65 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.692328 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 149.540000 0.000000 149.920000 0.900000 ;
    END
  END instr_rdata_i[25]
  PIN instr_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4854 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.857 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6255 LAYER met2  ;
    ANTENNAMAXAREACAR 23.4687 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 105.411 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.460000 0.000000 150.840000 0.900000 ;
    END
  END instr_rdata_i[24]
  PIN instr_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1914 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.515 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6255 LAYER met2  ;
    ANTENNAMAXAREACAR 22.6453 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 108.854 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 151.840000 0.000000 152.220000 0.900000 ;
    END
  END instr_rdata_i[23]
  PIN instr_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.2908 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.304 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6255 LAYER met2  ;
    ANTENNAMAXAREACAR 21.6141 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 94.3531 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 153.220000 0.000000 153.600000 0.900000 ;
    END
  END instr_rdata_i[22]
  PIN instr_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6121 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6255 LAYER met4  ;
    ANTENNAMAXAREACAR 21.6409 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 100.86 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.789346 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 154.600000 0.000000 154.980000 0.900000 ;
    END
  END instr_rdata_i[21]
  PIN instr_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7598 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.638 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.0858 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.928 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6255 LAYER met3  ;
    ANTENNAMAXAREACAR 34.8426 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 168.363 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.413796 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 155.520000 0.000000 155.900000 0.900000 ;
    END
  END instr_rdata_i[20]
  PIN instr_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7211 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.9725 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 19.2438 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 89.996 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.460202 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.1888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.144 LAYER met3  ;
    ANTENNAGATEAREA 0.6255 LAYER met3  ;
    ANTENNAMAXAREACAR 22.7431 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 109.411 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.692328 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 156.900000 0.000000 157.280000 0.900000 ;
    END
  END instr_rdata_i[19]
  PIN instr_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2533 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.1055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.5576 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 41.248 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6255 LAYER met4  ;
    ANTENNAMAXAREACAR 64.9252 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 326.264 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32725 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 158.280000 0.000000 158.660000 0.900000 ;
    END
  END instr_rdata_i[18]
  PIN instr_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4941 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 127.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.0697 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.504 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6255 LAYER met4  ;
    ANTENNAMAXAREACAR 35.2188 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 184.549 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.798148 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 159.660000 0.000000 160.040000 0.900000 ;
    END
  END instr_rdata_i[17]
  PIN instr_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7697 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.8265 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4995 LAYER met2  ;
    ANTENNAMAXAREACAR 28.5462 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 127.949 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.845159 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAGATEAREA 0.4995 LAYER met3  ;
    ANTENNAMAXAREACAR 29.0846 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 131.617 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.92524 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.6082 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 31.792 LAYER met4  ;
    ANTENNAGATEAREA 0.6255 LAYER met4  ;
    ANTENNAMAXAREACAR 38.0506 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 182.443 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 161.040000 0.000000 161.420000 0.900000 ;
    END
  END instr_rdata_i[16]
  PIN instr_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.9766 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.496 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 73.0702 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 351.258 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.9619 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.592 LAYER met3  ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 76.8873 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 373.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.884127 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.936 LAYER met4  ;
    ANTENNAGATEAREA 0.6255 LAYER met4  ;
    ANTENNAMAXAREACAR 79.1252 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 386.136 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.884127 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 161.960000 0.000000 162.340000 0.900000 ;
    END
  END instr_rdata_i[15]
  PIN instr_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.0686 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.655 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6255 LAYER met2  ;
    ANTENNAMAXAREACAR 24.4046 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 109.044 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 163.340000 0.000000 163.720000 0.900000 ;
    END
  END instr_rdata_i[14]
  PIN instr_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0997 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.593 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 110.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.1515 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.744 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6255 LAYER met4  ;
    ANTENNAMAXAREACAR 40.4905 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 202.138 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.85635 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 164.720000 0.000000 165.100000 0.900000 ;
    END
  END instr_rdata_i[13]
  PIN instr_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.7546 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.859 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6255 LAYER met2  ;
    ANTENNAMAXAREACAR 21.0286 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 92.66 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 166.100000 0.000000 166.480000 0.900000 ;
    END
  END instr_rdata_i[12]
  PIN instr_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3413 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.18348 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.432 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 34.4658 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 166.634 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.622127 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.3278 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.552 LAYER met4  ;
    ANTENNAGATEAREA 0.6255 LAYER met4  ;
    ANTENNAMAXAREACAR 41.3847 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 204.287 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 167.020000 0.000000 167.400000 0.900000 ;
    END
  END instr_rdata_i[11]
  PIN instr_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.732 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.09 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6255 LAYER met2  ;
    ANTENNAMAXAREACAR 24.479 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 110.14 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 168.400000 0.000000 168.780000 0.900000 ;
    END
  END instr_rdata_i[10]
  PIN instr_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4522 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.573 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6255 LAYER met2  ;
    ANTENNAMAXAREACAR 22.3179 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 98.6105 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 169.780000 0.000000 170.160000 0.900000 ;
    END
  END instr_rdata_i[9]
  PIN instr_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3122 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.767 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 22.7137 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 107.404 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.7696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.712 LAYER met3  ;
    ANTENNAGATEAREA 0.6255 LAYER met3  ;
    ANTENNAMAXAREACAR 46.3262 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 234.841 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 171.160000 0.000000 171.540000 0.900000 ;
    END
  END instr_rdata_i[8]
  PIN instr_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.402 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.3746 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.272 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6255 LAYER met4  ;
    ANTENNAMAXAREACAR 55.7339 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 280.705 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.864647 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 172.540000 0.000000 172.920000 0.900000 ;
    END
  END instr_rdata_i[7]
  PIN instr_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5629 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.096 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.7746 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 71.424 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6255 LAYER met4  ;
    ANTENNAMAXAREACAR 82.2202 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 432.282 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.36032 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 173.460000 0.000000 173.840000 0.900000 ;
    END
  END instr_rdata_i[6]
  PIN instr_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8213 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.5915 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 52.9782 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 248.925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 61.0813 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 295.845 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER met4  ;
    ANTENNAGATEAREA 0.6255 LAYER met4  ;
    ANTENNAMAXAREACAR 64.4895 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 314.774 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 174.840000 0.000000 175.220000 0.900000 ;
    END
  END instr_rdata_i[5]
  PIN instr_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7495 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.1345 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 28.3491 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 129.083 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.515032 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.2419 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.752 LAYER met3  ;
    ANTENNAGATEAREA 0.4995 LAYER met3  ;
    ANTENNAMAXAREACAR 58.8634 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 292.75 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.805477 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.7898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.016 LAYER met4  ;
    ANTENNAGATEAREA 0.6255 LAYER met4  ;
    ANTENNAMAXAREACAR 61.7248 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 308.763 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 176.220000 0.000000 176.600000 0.900000 ;
    END
  END instr_rdata_i[4]
  PIN instr_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2573 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.7815 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 13.8339 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 64.0025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.515032 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 14.5057 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 68.8432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.622127 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.3954 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.52 LAYER met4  ;
    ANTENNAGATEAREA 0.6255 LAYER met4  ;
    ANTENNAMAXAREACAR 24.7302 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 125.63 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 177.600000 0.000000 177.980000 0.900000 ;
    END
  END instr_rdata_i[3]
  PIN instr_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.2446 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.761 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6255 LAYER met2  ;
    ANTENNAMAXAREACAR 30.886 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 141.812 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 178.520000 0.000000 178.900000 0.900000 ;
    END
  END instr_rdata_i[2]
  PIN instr_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.6166 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.513 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6255 LAYER met2  ;
    ANTENNAMAXAREACAR 23.3542 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 103.981 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 179.900000 0.000000 180.280000 0.900000 ;
    END
  END instr_rdata_i[1]
  PIN instr_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.1806 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.989 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6255 LAYER met2  ;
    ANTENNAMAXAREACAR 34.7435 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 160.377 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 181.280000 0.000000 181.660000 0.900000 ;
    END
  END instr_rdata_i[0]
  PIN instr_rdata_intg_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.660000 0.000000 183.040000 0.900000 ;
    END
  END instr_rdata_intg_i[6]
  PIN instr_rdata_intg_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.040000 0.000000 184.420000 0.900000 ;
    END
  END instr_rdata_intg_i[5]
  PIN instr_rdata_intg_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.960000 0.000000 185.340000 0.900000 ;
    END
  END instr_rdata_intg_i[4]
  PIN instr_rdata_intg_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.340000 0.000000 186.720000 0.900000 ;
    END
  END instr_rdata_intg_i[3]
  PIN instr_rdata_intg_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.720000 0.000000 188.100000 0.900000 ;
    END
  END instr_rdata_intg_i[2]
  PIN instr_rdata_intg_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.100000 0.000000 189.480000 0.900000 ;
    END
  END instr_rdata_intg_i[1]
  PIN instr_rdata_intg_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.480000 0.000000 190.860000 0.900000 ;
    END
  END instr_rdata_intg_i[0]
  PIN instr_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.344 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 15.6671 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 73.623 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 191.400000 0.000000 191.780000 0.900000 ;
    END
  END instr_err_i
  PIN data_req_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4168 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.858 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 192.780000 0.000000 193.160000 0.900000 ;
    END
  END data_req_o
  PIN data_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.5706 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.746 LAYER met4  ;
    ANTENNAMAXAREACAR 19.639 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 86.0307 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.898187 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 194.160000 0.000000 194.540000 0.900000 ;
    END
  END data_gnt_i
  PIN data_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.9386 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 91.28 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 41.7915 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 218.803 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.555253 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 195.540000 0.000000 195.920000 0.900000 ;
    END
  END data_rvalid_i
  PIN data_we_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7626 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.587 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 196.460000 0.000000 196.840000 0.900000 ;
    END
  END data_we_o
  PIN data_be_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6986 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.267 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 197.840000 0.000000 198.220000 0.900000 ;
    END
  END data_be_o[3]
  PIN data_be_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.7538 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 53.543 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 199.220000 0.000000 199.600000 0.900000 ;
    END
  END data_be_o[2]
  PIN data_be_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.058 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 200.600000 0.000000 200.980000 0.900000 ;
    END
  END data_be_o[1]
  PIN data_be_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.498 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.264 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 201.980000 0.000000 202.360000 0.900000 ;
    END
  END data_be_o[0]
  PIN data_addr_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.5522 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 72.653 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 202.900000 0.000000 203.280000 0.900000 ;
    END
  END data_addr_o[31]
  PIN data_addr_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9971 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.8245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.1118 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 102.4 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 204.280000 0.000000 204.660000 0.900000 ;
    END
  END data_addr_o[30]
  PIN data_addr_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7362 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 205.660000 0.000000 206.040000 0.900000 ;
    END
  END data_addr_o[29]
  PIN data_addr_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.039 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.087 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 207.040000 0.000000 207.420000 0.900000 ;
    END
  END data_addr_o[28]
  PIN data_addr_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0318 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.933 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 207.960000 0.000000 208.340000 0.900000 ;
    END
  END data_addr_o[27]
  PIN data_addr_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6582 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.183 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.340000 0.000000 209.720000 0.900000 ;
    END
  END data_addr_o[26]
  PIN data_addr_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.127 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 210.720000 0.000000 211.100000 0.900000 ;
    END
  END data_addr_o[25]
  PIN data_addr_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.7116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.44 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 212.100000 0.000000 212.480000 0.900000 ;
    END
  END data_addr_o[24]
  PIN data_addr_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.4842 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.313 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 213.480000 0.000000 213.860000 0.900000 ;
    END
  END data_addr_o[23]
  PIN data_addr_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.079 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 214.400000 0.000000 214.780000 0.900000 ;
    END
  END data_addr_o[22]
  PIN data_addr_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.2918 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.351 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 215.780000 0.000000 216.160000 0.900000 ;
    END
  END data_addr_o[21]
  PIN data_addr_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.465 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.217 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 217.160000 0.000000 217.540000 0.900000 ;
    END
  END data_addr_o[20]
  PIN data_addr_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.306 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.304 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 218.540000 0.000000 218.920000 0.900000 ;
    END
  END data_addr_o[19]
  PIN data_addr_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.9586 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.685 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 219.460000 0.000000 219.840000 0.900000 ;
    END
  END data_addr_o[18]
  PIN data_addr_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.135 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.567 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 220.840000 0.000000 221.220000 0.900000 ;
    END
  END data_addr_o[17]
  PIN data_addr_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6246 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.015 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 222.220000 0.000000 222.600000 0.900000 ;
    END
  END data_addr_o[16]
  PIN data_addr_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9102 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.443 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 223.600000 0.000000 223.980000 0.900000 ;
    END
  END data_addr_o[15]
  PIN data_addr_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.8934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.359 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 224.980000 0.000000 225.360000 0.900000 ;
    END
  END data_addr_o[14]
  PIN data_addr_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9578 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.681 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 225.900000 0.000000 226.280000 0.900000 ;
    END
  END data_addr_o[13]
  PIN data_addr_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.435 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 227.280000 0.000000 227.660000 0.900000 ;
    END
  END data_addr_o[12]
  PIN data_addr_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.7733 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.7585 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 228.660000 0.000000 229.040000 0.900000 ;
    END
  END data_addr_o[11]
  PIN data_addr_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.672 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.134 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 230.040000 0.000000 230.420000 0.900000 ;
    END
  END data_addr_o[10]
  PIN data_addr_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.5246 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.397 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 230.960000 0.000000 231.340000 0.900000 ;
    END
  END data_addr_o[9]
  PIN data_addr_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.6565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.0878 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 86.272 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 232.340000 0.000000 232.720000 0.900000 ;
    END
  END data_addr_o[8]
  PIN data_addr_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2374 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.843 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 233.720000 0.000000 234.100000 0.900000 ;
    END
  END data_addr_o[7]
  PIN data_addr_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0143 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.6978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 84.192 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 235.100000 0.000000 235.480000 0.900000 ;
    END
  END data_addr_o[6]
  PIN data_addr_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0143 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.8438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.304 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 236.480000 0.000000 236.860000 0.900000 ;
    END
  END data_addr_o[5]
  PIN data_addr_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.849 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.4818 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 131.04 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 237.400000 0.000000 237.780000 0.900000 ;
    END
  END data_addr_o[4]
  PIN data_addr_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2966 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.375 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 238.780000 0.000000 239.160000 0.900000 ;
    END
  END data_addr_o[3]
  PIN data_addr_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.3188 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 103.504 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 240.160000 0.000000 240.540000 0.900000 ;
    END
  END data_addr_o[2]
  PIN data_addr_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3722 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.753 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 241.540000 0.000000 241.920000 0.900000 ;
    END
  END data_addr_o[1]
  PIN data_addr_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0787 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.2298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.696 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 242.460000 0.000000 242.840000 0.900000 ;
    END
  END data_addr_o[0]
  PIN data_wdata_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4058 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.921 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 243.840000 0.000000 244.220000 0.900000 ;
    END
  END data_wdata_o[31]
  PIN data_wdata_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.6934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.359 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 245.220000 0.000000 245.600000 0.900000 ;
    END
  END data_wdata_o[30]
  PIN data_wdata_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5558 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.553 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 246.600000 0.000000 246.980000 0.900000 ;
    END
  END data_wdata_o[29]
  PIN data_wdata_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4986 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.385 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 247.980000 0.000000 248.360000 0.900000 ;
    END
  END data_wdata_o[28]
  PIN data_wdata_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.837 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 248.900000 0.000000 249.280000 0.900000 ;
    END
  END data_wdata_o[27]
  PIN data_wdata_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.0002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.775 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 250.280000 0.000000 250.660000 0.900000 ;
    END
  END data_wdata_o[26]
  PIN data_wdata_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.5368 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 78 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 251.660000 0.000000 252.040000 0.900000 ;
    END
  END data_wdata_o[25]
  PIN data_wdata_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.5718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.633 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 253.040000 0.000000 253.420000 0.900000 ;
    END
  END data_wdata_o[24]
  PIN data_wdata_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9914 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.849 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 254.420000 0.000000 254.800000 0.900000 ;
    END
  END data_wdata_o[23]
  PIN data_wdata_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1606 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.577 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 255.340000 0.000000 255.720000 0.900000 ;
    END
  END data_wdata_o[22]
  PIN data_wdata_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0143 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.2618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 135.2 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 256.720000 0.000000 257.100000 0.900000 ;
    END
  END data_wdata_o[21]
  PIN data_wdata_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8626 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.205 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 258.100000 0.000000 258.480000 0.900000 ;
    END
  END data_wdata_o[20]
  PIN data_wdata_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.935 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 259.480000 0.000000 259.860000 0.900000 ;
    END
  END data_wdata_o[19]
  PIN data_wdata_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0143 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.1598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.656 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 260.400000 0.000000 260.780000 0.900000 ;
    END
  END data_wdata_o[18]
  PIN data_wdata_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1773 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.263 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.9048 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 85.296 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 261.780000 0.000000 262.160000 0.900000 ;
    END
  END data_wdata_o[17]
  PIN data_wdata_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9537 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.93 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.76 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.6958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 62.848 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 263.160000 0.000000 263.540000 0.900000 ;
    END
  END data_wdata_o[16]
  PIN data_wdata_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0143 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.8198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 90.176 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 264.540000 0.000000 264.920000 0.900000 ;
    END
  END data_wdata_o[15]
  PIN data_wdata_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.2838 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 97.984 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 265.920000 0.000000 266.300000 0.900000 ;
    END
  END data_wdata_o[14]
  PIN data_wdata_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.5634 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.709 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 266.840000 0.000000 267.220000 0.900000 ;
    END
  END data_wdata_o[13]
  PIN data_wdata_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4413 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.7918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 31.36 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 268.220000 0.000000 268.600000 0.900000 ;
    END
  END data_wdata_o[12]
  PIN data_wdata_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.5798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 152.896 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 269.600000 0.000000 269.980000 0.900000 ;
    END
  END data_wdata_o[11]
  PIN data_wdata_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6034 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.791 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 270.980000 0.000000 271.360000 0.900000 ;
    END
  END data_wdata_o[10]
  PIN data_wdata_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.354 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.1468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 59.92 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 271.900000 0.000000 272.280000 0.900000 ;
    END
  END data_wdata_o[9]
  PIN data_wdata_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6034 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.791 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 273.280000 0.000000 273.660000 0.900000 ;
    END
  END data_wdata_o[8]
  PIN data_wdata_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6244 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.896 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 274.660000 0.000000 275.040000 0.900000 ;
    END
  END data_wdata_o[7]
  PIN data_wdata_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.0158 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 101.888 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 276.040000 0.000000 276.420000 0.900000 ;
    END
  END data_wdata_o[6]
  PIN data_wdata_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.63 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 277.420000 0.000000 277.800000 0.900000 ;
    END
  END data_wdata_o[5]
  PIN data_wdata_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5057 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.0178 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 139.232 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 278.340000 0.000000 278.720000 0.900000 ;
    END
  END data_wdata_o[4]
  PIN data_wdata_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5451 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.2488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 156.464 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 279.720000 0.000000 280.100000 0.900000 ;
    END
  END data_wdata_o[3]
  PIN data_wdata_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9264 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 281.100000 0.000000 281.480000 0.900000 ;
    END
  END data_wdata_o[2]
  PIN data_wdata_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0318 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.933 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 282.480000 0.000000 282.860000 0.900000 ;
    END
  END data_wdata_o[1]
  PIN data_wdata_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7054 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.419 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 283.400000 0.000000 283.780000 0.900000 ;
    END
  END data_wdata_o[0]
  PIN data_wdata_intg_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.44 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.082 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 284.780000 0.000000 285.160000 0.900000 ;
    END
  END data_wdata_intg_o[6]
  PIN data_wdata_intg_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.41 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.942 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 286.160000 0.000000 286.540000 0.900000 ;
    END
  END data_wdata_intg_o[5]
  PIN data_wdata_intg_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.563 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.707 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 287.540000 0.000000 287.920000 0.900000 ;
    END
  END data_wdata_intg_o[4]
  PIN data_wdata_intg_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6202 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.875 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 288.920000 0.000000 289.300000 0.900000 ;
    END
  END data_wdata_intg_o[3]
  PIN data_wdata_intg_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1674 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.729 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 289.840000 0.000000 290.220000 0.900000 ;
    END
  END data_wdata_intg_o[2]
  PIN data_wdata_intg_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3174 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.361 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 291.220000 0.000000 291.600000 0.900000 ;
    END
  END data_wdata_intg_o[1]
  PIN data_wdata_intg_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.103 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.407 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 292.600000 0.000000 292.980000 0.900000 ;
    END
  END data_wdata_intg_o[0]
  PIN data_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0143 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.6784 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 143.696 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 60.0573 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 317.599 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.35025 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 293.980000 0.000000 294.360000 0.900000 ;
    END
  END data_rdata_i[31]
  PIN data_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4775 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.0519 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 130.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 93.8349 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 485.132 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.36032 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 294.900000 0.000000 295.280000 0.900000 ;
    END
  END data_rdata_i[30]
  PIN data_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.266 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.392 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 105.296 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 46.8718 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 234.62 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 296.280000 0.000000 296.660000 0.900000 ;
    END
  END data_rdata_i[29]
  PIN data_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1431 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 60.0156 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 321.024 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 85.2659 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 433.94 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.771453 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 297.660000 0.000000 298.040000 0.900000 ;
    END
  END data_rdata_i[28]
  PIN data_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3935 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.8065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 53.1021 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 285.088 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 84.5845 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 428.319 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.536761 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 299.040000 0.000000 299.420000 0.900000 ;
    END
  END data_rdata_i[27]
  PIN data_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9539 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.059 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.2413 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 141.36 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 65.9618 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 346.016 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.832492 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 300.420000 0.000000 300.800000 0.900000 ;
    END
  END data_rdata_i[26]
  PIN data_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0787 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 23.1366 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 124.336 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 102.266 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 523.68 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.854221 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 301.340000 0.000000 301.720000 0.900000 ;
    END
  END data_rdata_i[25]
  PIN data_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6525 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.485 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.8473 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 80.592 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 28.1335 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 151.207 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 302.720000 0.000000 303.100000 0.900000 ;
    END
  END data_rdata_i[24]
  PIN data_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.0586 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 45.4063 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 230.621 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.771453 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 304.100000 0.000000 304.480000 0.900000 ;
    END
  END data_rdata_i[23]
  PIN data_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0716 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.916 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 13.601 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 50.2542 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 305.480000 0.000000 305.860000 0.900000 ;
    END
  END data_rdata_i[22]
  PIN data_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8263 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.9705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.9626 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.408 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 76.5052 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 387.162 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.854221 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 306.860000 0.000000 307.240000 0.900000 ;
    END
  END data_rdata_i[21]
  PIN data_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6555 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 55.1454 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 295.52 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 77.7383 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 393.003 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.678621 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 307.780000 0.000000 308.160000 0.900000 ;
    END
  END data_rdata_i[20]
  PIN data_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6975 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.4684 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 222.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 67.6212 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 353.983 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.518405 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 309.160000 0.000000 309.540000 0.900000 ;
    END
  END data_rdata_i[19]
  PIN data_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2821 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.931 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.5044 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 62.768 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 45.4493 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 240.203 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.692525 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 310.540000 0.000000 310.920000 0.900000 ;
    END
  END data_rdata_i[18]
  PIN data_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 44.9226 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 240.528 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 74.8826 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 393.372 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.771453 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 311.920000 0.000000 312.300000 0.900000 ;
    END
  END data_rdata_i[17]
  PIN data_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3559 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.2754 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 66.88 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 47.2833 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 249.713 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.854221 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 312.840000 0.000000 313.220000 0.900000 ;
    END
  END data_rdata_i[16]
  PIN data_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.936 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 44.4505 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 209.185 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.678621 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 314.220000 0.000000 314.600000 0.900000 ;
    END
  END data_rdata_i[15]
  PIN data_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.0545 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 14.738 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 68.897 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.0848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.256 LAYER met3  ;
    ANTENNAGATEAREA 0.8685 LAYER met3  ;
    ANTENNAMAXAREACAR 15.987 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 76.1002 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.65092 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 315.600000 0.000000 315.980000 0.900000 ;
    END
  END data_rdata_i[14]
  PIN data_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1431 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.4538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 120.672 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 79.9894 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 403.173 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.729222 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4  ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 84.7618 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 429.168 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.729222 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 316.980000 0.000000 317.360000 0.900000 ;
    END
  END data_rdata_i[13]
  PIN data_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2041 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.7858 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 159.328 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met3  ;
    ANTENNAMAXAREACAR 49.0863 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 239.034 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.453993 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 318.360000 0.000000 318.740000 0.900000 ;
    END
  END data_rdata_i[12]
  PIN data_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3233 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.849 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.1644 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 50.288 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 93.7887 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 496.912 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.854141 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 319.280000 0.000000 319.660000 0.900000 ;
    END
  END data_rdata_i[11]
  PIN data_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.86 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 29.9769 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 130.754 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.515032 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.6028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.352 LAYER met3  ;
    ANTENNAGATEAREA 0.8685 LAYER met3  ;
    ANTENNAMAXAREACAR 32.9737 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 147.279 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.515032 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 320.660000 0.000000 321.040000 0.900000 ;
    END
  END data_rdata_i[10]
  PIN data_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7982 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.539 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 16.6198 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 64.8006 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 322.040000 0.000000 322.420000 0.900000 ;
    END
  END data_rdata_i[9]
  PIN data_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.2161 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.3395 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 17.986 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 70.959 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.472349 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.7748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAGATEAREA 0.8685 LAYER met3  ;
    ANTENNAMAXAREACAR 20.0295 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 82.3994 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.472349 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 323.420000 0.000000 323.800000 0.900000 ;
    END
  END data_rdata_i[8]
  PIN data_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.395 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.4018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 45.28 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 32.3771 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 149.056 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.715332 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 324.340000 0.000000 324.720000 0.900000 ;
    END
  END data_rdata_i[7]
  PIN data_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5556 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.552 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 14.801 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 55.8632 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 325.720000 0.000000 326.100000 0.900000 ;
    END
  END data_rdata_i[6]
  PIN data_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3793 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2413 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1046 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 23.0346 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 102.593 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.536761 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 327.100000 0.000000 327.480000 0.900000 ;
    END
  END data_rdata_i[5]
  PIN data_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7512 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.52 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 25.0549 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 106.259 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 328.480000 0.000000 328.860000 0.900000 ;
    END
  END data_rdata_i[4]
  PIN data_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9045 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.1208 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 38.448 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 23.7807 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 111.904 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.789809 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 329.860000 0.000000 330.240000 0.900000 ;
    END
  END data_rdata_i[3]
  PIN data_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2653 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.58 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 147.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.5218 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 23.1653 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 103.913 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.789809 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 330.780000 0.000000 331.160000 0.900000 ;
    END
  END data_rdata_i[2]
  PIN data_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1978 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.655 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 15.247 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 57.9195 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 332.160000 0.000000 332.540000 0.900000 ;
    END
  END data_rdata_i[1]
  PIN data_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2368 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 15.3098 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 58.0435 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 333.540000 0.000000 333.920000 0.900000 ;
    END
  END data_rdata_i[0]
  PIN data_rdata_intg_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.920000 0.000000 335.300000 0.900000 ;
    END
  END data_rdata_intg_i[6]
  PIN data_rdata_intg_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.840000 0.000000 336.220000 0.900000 ;
    END
  END data_rdata_intg_i[5]
  PIN data_rdata_intg_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.220000 0.000000 337.600000 0.900000 ;
    END
  END data_rdata_intg_i[4]
  PIN data_rdata_intg_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.600000 0.000000 338.980000 0.900000 ;
    END
  END data_rdata_intg_i[3]
  PIN data_rdata_intg_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.980000 0.000000 340.360000 0.900000 ;
    END
  END data_rdata_intg_i[2]
  PIN data_rdata_intg_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.360000 0.000000 341.740000 0.900000 ;
    END
  END data_rdata_intg_i[1]
  PIN data_rdata_intg_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.280000 0.000000 342.660000 0.900000 ;
    END
  END data_rdata_intg_i[0]
  PIN data_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2503 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.9725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.4758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 43.7206 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 220.939 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.536761 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 343.660000 0.000000 344.040000 0.900000 ;
    END
  END data_err_i
  PIN eFPGA_operand_a_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 24.3264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 129.736 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 9.840000 550.160000 10.220000 ;
    END
  END eFPGA_operand_a_o[31]
  PIN eFPGA_operand_a_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.1466 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 171.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.3908 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 55.888 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 12.890000 550.160000 13.270000 ;
    END
  END eFPGA_operand_a_o[30]
  PIN eFPGA_operand_a_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.8074 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.968 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 16.550000 550.160000 16.930000 ;
    END
  END eFPGA_operand_a_o[29]
  PIN eFPGA_operand_a_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.3664 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 158.032 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 19.600000 550.160000 19.980000 ;
    END
  END eFPGA_operand_a_o[28]
  PIN eFPGA_operand_a_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3346 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.5298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 115.296 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 23.260000 550.160000 23.640000 ;
    END
  END eFPGA_operand_a_o[27]
  PIN eFPGA_operand_a_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3476 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.9238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 176.064 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 26.920000 550.160000 27.300000 ;
    END
  END eFPGA_operand_a_o[26]
  PIN eFPGA_operand_a_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2456 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.0796 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 188.032 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 29.970000 550.160000 30.350000 ;
    END
  END eFPGA_operand_a_o[25]
  PIN eFPGA_operand_a_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7896 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.3956 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 168.384 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 33.630000 550.160000 34.010000 ;
    END
  END eFPGA_operand_a_o[24]
  PIN eFPGA_operand_a_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.7704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.104 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 37.290000 550.160000 37.670000 ;
    END
  END eFPGA_operand_a_o[23]
  PIN eFPGA_operand_a_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.6022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 142.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 40.340000 550.160000 40.720000 ;
    END
  END eFPGA_operand_a_o[22]
  PIN eFPGA_operand_a_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.3424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.488 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 44.000000 550.160000 44.380000 ;
    END
  END eFPGA_operand_a_o[21]
  PIN eFPGA_operand_a_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 47.660000 550.160000 48.040000 ;
    END
  END eFPGA_operand_a_o[20]
  PIN eFPGA_operand_a_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5594 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.312 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 50.710000 550.160000 51.090000 ;
    END
  END eFPGA_operand_a_o[19]
  PIN eFPGA_operand_a_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.7564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.696 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 54.370000 550.160000 54.750000 ;
    END
  END eFPGA_operand_a_o[18]
  PIN eFPGA_operand_a_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 58.030000 550.160000 58.410000 ;
    END
  END eFPGA_operand_a_o[17]
  PIN eFPGA_operand_a_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.1452 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 61.080000 550.160000 61.460000 ;
    END
  END eFPGA_operand_a_o[16]
  PIN eFPGA_operand_a_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.5198 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 120.576 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 64.740000 550.160000 65.120000 ;
    END
  END eFPGA_operand_a_o[15]
  PIN eFPGA_operand_a_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.2852 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 119.32 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 68.400000 550.160000 68.780000 ;
    END
  END eFPGA_operand_a_o[14]
  PIN eFPGA_operand_a_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.1704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.904 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 71.450000 550.160000 71.830000 ;
    END
  END eFPGA_operand_a_o[13]
  PIN eFPGA_operand_a_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.1472 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 118.584 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 75.110000 550.160000 75.490000 ;
    END
  END eFPGA_operand_a_o[12]
  PIN eFPGA_operand_a_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.5844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.112 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 78.770000 550.160000 79.150000 ;
    END
  END eFPGA_operand_a_o[11]
  PIN eFPGA_operand_a_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.5954 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 81.820000 550.160000 82.200000 ;
    END
  END eFPGA_operand_a_o[10]
  PIN eFPGA_operand_a_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6864 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.656 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 85.480000 550.160000 85.860000 ;
    END
  END eFPGA_operand_a_o[9]
  PIN eFPGA_operand_a_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 89.140000 550.160000 89.520000 ;
    END
  END eFPGA_operand_a_o[8]
  PIN eFPGA_operand_a_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 92.190000 550.160000 92.570000 ;
    END
  END eFPGA_operand_a_o[7]
  PIN eFPGA_operand_a_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.1844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.312 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 95.850000 550.160000 96.230000 ;
    END
  END eFPGA_operand_a_o[6]
  PIN eFPGA_operand_a_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 99.510000 550.160000 99.890000 ;
    END
  END eFPGA_operand_a_o[5]
  PIN eFPGA_operand_a_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.5024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.008 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 102.560000 550.160000 102.940000 ;
    END
  END eFPGA_operand_a_o[4]
  PIN eFPGA_operand_a_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 106.220000 550.160000 106.600000 ;
    END
  END eFPGA_operand_a_o[3]
  PIN eFPGA_operand_a_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.4124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.528 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 109.270000 550.160000 109.650000 ;
    END
  END eFPGA_operand_a_o[2]
  PIN eFPGA_operand_a_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 23.3802 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125.16 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 112.930000 550.160000 113.310000 ;
    END
  END eFPGA_operand_a_o[1]
  PIN eFPGA_operand_a_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7616 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.4138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 205.344 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 116.590000 550.160000 116.970000 ;
    END
  END eFPGA_operand_a_o[0]
  PIN eFPGA_operand_b_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.4464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.376 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 119.640000 550.160000 120.020000 ;
    END
  END eFPGA_operand_b_o[31]
  PIN eFPGA_operand_b_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 123.300000 550.160000 123.680000 ;
    END
  END eFPGA_operand_b_o[30]
  PIN eFPGA_operand_b_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 32.3724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 172.648 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 126.960000 550.160000 127.340000 ;
    END
  END eFPGA_operand_b_o[29]
  PIN eFPGA_operand_b_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9076 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.936 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 130.010000 550.160000 130.390000 ;
    END
  END eFPGA_operand_b_o[28]
  PIN eFPGA_operand_b_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.2964 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.576 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 133.670000 550.160000 134.050000 ;
    END
  END eFPGA_operand_b_o[27]
  PIN eFPGA_operand_b_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.2264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.536 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 137.330000 550.160000 137.710000 ;
    END
  END eFPGA_operand_b_o[26]
  PIN eFPGA_operand_b_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.6196 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 140.380000 550.160000 140.760000 ;
    END
  END eFPGA_operand_b_o[25]
  PIN eFPGA_operand_b_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.2914 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 92.216 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 144.040000 550.160000 144.420000 ;
    END
  END eFPGA_operand_b_o[24]
  PIN eFPGA_operand_b_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.1364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.056 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 147.700000 550.160000 148.080000 ;
    END
  END eFPGA_operand_b_o[23]
  PIN eFPGA_operand_b_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 150.750000 550.160000 151.130000 ;
    END
  END eFPGA_operand_b_o[22]
  PIN eFPGA_operand_b_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 154.410000 550.160000 154.790000 ;
    END
  END eFPGA_operand_b_o[21]
  PIN eFPGA_operand_b_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 158.070000 550.160000 158.450000 ;
    END
  END eFPGA_operand_b_o[20]
  PIN eFPGA_operand_b_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.3174 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 161.120000 550.160000 161.500000 ;
    END
  END eFPGA_operand_b_o[19]
  PIN eFPGA_operand_b_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.2754 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.464 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 164.780000 550.160000 165.160000 ;
    END
  END eFPGA_operand_b_o[18]
  PIN eFPGA_operand_b_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.5504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.264 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 168.440000 550.160000 168.820000 ;
    END
  END eFPGA_operand_b_o[17]
  PIN eFPGA_operand_b_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 171.490000 550.160000 171.870000 ;
    END
  END eFPGA_operand_b_o[16]
  PIN eFPGA_operand_b_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.1634 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 118.2 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 175.150000 550.160000 175.530000 ;
    END
  END eFPGA_operand_b_o[15]
  PIN eFPGA_operand_b_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 178.810000 550.160000 179.190000 ;
    END
  END eFPGA_operand_b_o[14]
  PIN eFPGA_operand_b_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.0046 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 176.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 181.860000 550.160000 182.240000 ;
    END
  END eFPGA_operand_b_o[13]
  PIN eFPGA_operand_b_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4846 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.0806 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.704 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 185.520000 550.160000 185.900000 ;
    END
  END eFPGA_operand_b_o[12]
  PIN eFPGA_operand_b_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 189.180000 550.160000 189.560000 ;
    END
  END eFPGA_operand_b_o[11]
  PIN eFPGA_operand_b_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.8492 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 106.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 192.230000 550.160000 192.610000 ;
    END
  END eFPGA_operand_b_o[10]
  PIN eFPGA_operand_b_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.2804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.824 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 195.890000 550.160000 196.270000 ;
    END
  END eFPGA_operand_b_o[9]
  PIN eFPGA_operand_b_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.1494 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 112.792 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 199.550000 550.160000 199.930000 ;
    END
  END eFPGA_operand_b_o[8]
  PIN eFPGA_operand_b_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.9614 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 106.456 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 202.600000 550.160000 202.980000 ;
    END
  END eFPGA_operand_b_o[7]
  PIN eFPGA_operand_b_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.1514 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 134.136 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 206.260000 550.160000 206.640000 ;
    END
  END eFPGA_operand_b_o[6]
  PIN eFPGA_operand_b_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.9284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 209.310000 550.160000 209.690000 ;
    END
  END eFPGA_operand_b_o[5]
  PIN eFPGA_operand_b_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.1206 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 212.970000 550.160000 213.350000 ;
    END
  END eFPGA_operand_b_o[4]
  PIN eFPGA_operand_b_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 216.630000 550.160000 217.010000 ;
    END
  END eFPGA_operand_b_o[3]
  PIN eFPGA_operand_b_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 219.680000 550.160000 220.060000 ;
    END
  END eFPGA_operand_b_o[2]
  PIN eFPGA_operand_b_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.5844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.112 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 223.340000 550.160000 223.720000 ;
    END
  END eFPGA_operand_b_o[1]
  PIN eFPGA_operand_b_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 227.000000 550.160000 227.380000 ;
    END
  END eFPGA_operand_b_o[0]
  PIN eFPGA_result_a_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.928 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 66.2917 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 342.642 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 230.050000 550.160000 230.430000 ;
    END
  END eFPGA_result_a_i[31]
  PIN eFPGA_result_a_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0132 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.536 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 17.5889 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 87.996 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 233.710000 550.160000 234.090000 ;
    END
  END eFPGA_result_a_i[30]
  PIN eFPGA_result_a_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 15.9119 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 76.0364 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 237.370000 550.160000 237.750000 ;
    END
  END eFPGA_result_a_i[29]
  PIN eFPGA_result_a_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 79.3956 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 391.208 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 240.420000 550.160000 240.800000 ;
    END
  END eFPGA_result_a_i[28]
  PIN eFPGA_result_a_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2664 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 82.4727 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 410.497 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 244.080000 550.160000 244.460000 ;
    END
  END eFPGA_result_a_i[27]
  PIN eFPGA_result_a_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9154 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.0008 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 53.808 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 45.3244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 238.873 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 247.740000 550.160000 248.120000 ;
    END
  END eFPGA_result_a_i[26]
  PIN eFPGA_result_a_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 11.3624 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 51.4707 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 250.790000 550.160000 251.170000 ;
    END
  END eFPGA_result_a_i[25]
  PIN eFPGA_result_a_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 11.1681 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 50.2303 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 254.450000 550.160000 254.830000 ;
    END
  END eFPGA_result_a_i[24]
  PIN eFPGA_result_a_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 82.097 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 405.063 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 258.110000 550.160000 258.490000 ;
    END
  END eFPGA_result_a_i[23]
  PIN eFPGA_result_a_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.27 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.376 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 15.5469 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 80.0444 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 261.160000 550.160000 261.540000 ;
    END
  END eFPGA_result_a_i[22]
  PIN eFPGA_result_a_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.472 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 83.6485 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 416.109 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 264.820000 550.160000 265.200000 ;
    END
  END eFPGA_result_a_i[21]
  PIN eFPGA_result_a_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8014 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.936 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 44.1455 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 218.562 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 268.480000 550.160000 268.860000 ;
    END
  END eFPGA_result_a_i[20]
  PIN eFPGA_result_a_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.28 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 85.1281 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 422.448 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 271.530000 550.160000 271.910000 ;
    END
  END eFPGA_result_a_i[19]
  PIN eFPGA_result_a_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.336 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 81.9701 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 405.915 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 275.190000 550.160000 275.570000 ;
    END
  END eFPGA_result_a_i[18]
  PIN eFPGA_result_a_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.92 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 12.1616 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 55.6081 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 278.850000 550.160000 279.230000 ;
    END
  END eFPGA_result_a_i[17]
  PIN eFPGA_result_a_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.3278 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.552 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 88.9568 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 451.863 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 281.900000 550.160000 282.280000 ;
    END
  END eFPGA_result_a_i[16]
  PIN eFPGA_result_a_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.64 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 64.4299 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 317.636 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 285.560000 550.160000 285.940000 ;
    END
  END eFPGA_result_a_i[15]
  PIN eFPGA_result_a_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4914 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.616 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 83.3374 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 415.6 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 289.220000 550.160000 289.600000 ;
    END
  END eFPGA_result_a_i[14]
  PIN eFPGA_result_a_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.864 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 13.4145 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 63.1192 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 292.270000 550.160000 292.650000 ;
    END
  END eFPGA_result_a_i[13]
  PIN eFPGA_result_a_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6912 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.152 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 52.2747 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 266.497 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 295.930000 550.160000 296.310000 ;
    END
  END eFPGA_result_a_i[12]
  PIN eFPGA_result_a_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6184 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.96 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 26.596 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 130.533 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 299.590000 550.160000 299.970000 ;
    END
  END eFPGA_result_a_i[11]
  PIN eFPGA_result_a_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.376 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.608 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 44.6984 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 232.667 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 302.640000 550.160000 303.020000 ;
    END
  END eFPGA_result_a_i[10]
  PIN eFPGA_result_a_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 16.1844 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 85.0747 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 306.300000 550.160000 306.680000 ;
    END
  END eFPGA_result_a_i[9]
  PIN eFPGA_result_a_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.888 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 82.0461 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 408.202 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 309.350000 550.160000 309.730000 ;
    END
  END eFPGA_result_a_i[8]
  PIN eFPGA_result_a_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9088 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.92 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 53.8636 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 280.158 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 313.010000 550.160000 313.390000 ;
    END
  END eFPGA_result_a_i[7]
  PIN eFPGA_result_a_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5066 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.4368 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 34.8 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 84.6384 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 430.145 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 316.670000 550.160000 317.050000 ;
    END
  END eFPGA_result_a_i[6]
  PIN eFPGA_result_a_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.6938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.504 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 81.1564 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 410.832 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 319.720000 550.160000 320.100000 ;
    END
  END eFPGA_result_a_i[5]
  PIN eFPGA_result_a_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.904 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 79.1725 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 394.343 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 323.380000 550.160000 323.760000 ;
    END
  END eFPGA_result_a_i[4]
  PIN eFPGA_result_a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 28.5329 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 135.758 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 327.040000 550.160000 327.420000 ;
    END
  END eFPGA_result_a_i[3]
  PIN eFPGA_result_a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9624 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.128 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 12.4259 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 57.9111 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 330.090000 550.160000 330.470000 ;
    END
  END eFPGA_result_a_i[2]
  PIN eFPGA_result_a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.96 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 60.7539 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 298.327 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 333.750000 550.160000 334.130000 ;
    END
  END eFPGA_result_a_i[1]
  PIN eFPGA_result_a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7372 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.064 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 27.9943 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 139.293 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 337.410000 550.160000 337.790000 ;
    END
  END eFPGA_result_a_i[0]
  PIN eFPGA_result_b_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.616 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.888 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 56.5254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 285.778 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 340.460000 550.160000 340.840000 ;
    END
  END eFPGA_result_b_i[31]
  PIN eFPGA_result_b_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.92 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 81.0976 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 387.365 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 344.120000 550.160000 344.500000 ;
    END
  END eFPGA_result_b_i[30]
  PIN eFPGA_result_b_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 77.0524 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 381.27 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 347.780000 550.160000 348.160000 ;
    END
  END eFPGA_result_b_i[29]
  PIN eFPGA_result_b_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.888 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 65.8071 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 325.722 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 350.830000 550.160000 351.210000 ;
    END
  END eFPGA_result_b_i[28]
  PIN eFPGA_result_b_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3414 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.816 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 60.2825 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 299.016 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 354.490000 550.160000 354.870000 ;
    END
  END eFPGA_result_b_i[27]
  PIN eFPGA_result_b_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4914 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.616 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 55.9746 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 269.936 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 358.150000 550.160000 358.530000 ;
    END
  END eFPGA_result_b_i[26]
  PIN eFPGA_result_b_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.032 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 50.2238 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 243.373 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 361.200000 550.160000 361.580000 ;
    END
  END eFPGA_result_b_i[25]
  PIN eFPGA_result_b_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.096 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 72.5444 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 359.968 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 364.860000 550.160000 365.240000 ;
    END
  END eFPGA_result_b_i[24]
  PIN eFPGA_result_b_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.9414 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 76.3444 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 380.913 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 368.520000 550.160000 368.900000 ;
    END
  END eFPGA_result_b_i[23]
  PIN eFPGA_result_b_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.9884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 83.7095 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 420.508 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 371.570000 550.160000 371.950000 ;
    END
  END eFPGA_result_b_i[22]
  PIN eFPGA_result_b_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 59.7048 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 292.849 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 375.230000 550.160000 375.610000 ;
    END
  END eFPGA_result_b_i[21]
  PIN eFPGA_result_b_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7224 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.848 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 56.5079 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 273.214 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 378.890000 550.160000 379.270000 ;
    END
  END eFPGA_result_b_i[20]
  PIN eFPGA_result_b_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1134 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 63.6659 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 315.865 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 381.940000 550.160000 382.320000 ;
    END
  END eFPGA_result_b_i[19]
  PIN eFPGA_result_b_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 40.7603 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 187.905 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 385.600000 550.160000 385.980000 ;
    END
  END eFPGA_result_b_i[18]
  PIN eFPGA_result_b_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7044 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.752 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 66.2968 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 330.048 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 389.260000 550.160000 389.640000 ;
    END
  END eFPGA_result_b_i[17]
  PIN eFPGA_result_b_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.624 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 62.4984 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 309.008 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 392.310000 550.160000 392.690000 ;
    END
  END eFPGA_result_b_i[16]
  PIN eFPGA_result_b_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 35.527 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 161.738 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 395.970000 550.160000 396.350000 ;
    END
  END eFPGA_result_b_i[15]
  PIN eFPGA_result_b_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 32.854 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 145.135 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 399.020000 550.160000 399.400000 ;
    END
  END eFPGA_result_b_i[14]
  PIN eFPGA_result_b_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2964 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 61.0984 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 303 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 402.680000 550.160000 403.060000 ;
    END
  END eFPGA_result_b_i[13]
  PIN eFPGA_result_b_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.392 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 34.4857 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 155.437 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 406.340000 550.160000 406.720000 ;
    END
  END eFPGA_result_b_i[12]
  PIN eFPGA_result_b_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3894 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.072 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 59.8333 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 296.825 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 409.390000 550.160000 409.770000 ;
    END
  END eFPGA_result_b_i[11]
  PIN eFPGA_result_b_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.5384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 66.8762 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 334.627 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 413.050000 550.160000 413.430000 ;
    END
  END eFPGA_result_b_i[10]
  PIN eFPGA_result_b_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6544 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.152 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 57.019 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 280.881 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 416.710000 550.160000 417.090000 ;
    END
  END eFPGA_result_b_i[9]
  PIN eFPGA_result_b_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.9864 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.256 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 65.5937 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 327.206 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 419.760000 550.160000 420.140000 ;
    END
  END eFPGA_result_b_i[8]
  PIN eFPGA_result_b_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.392 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 31.8968 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 142.492 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 423.420000 550.160000 423.800000 ;
    END
  END eFPGA_result_b_i[7]
  PIN eFPGA_result_b_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 51.6413 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 254.317 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 427.080000 550.160000 427.460000 ;
    END
  END eFPGA_result_b_i[6]
  PIN eFPGA_result_b_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.16 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 53.6095 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 263.341 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 430.130000 550.160000 430.510000 ;
    END
  END eFPGA_result_b_i[5]
  PIN eFPGA_result_b_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.864 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 33.5873 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 151.675 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 433.790000 550.160000 434.170000 ;
    END
  END eFPGA_result_b_i[4]
  PIN eFPGA_result_b_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 50.0095 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 245.19 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 437.450000 550.160000 437.830000 ;
    END
  END eFPGA_result_b_i[3]
  PIN eFPGA_result_b_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.056 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 39.7238 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 190.794 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 440.500000 550.160000 440.880000 ;
    END
  END eFPGA_result_b_i[2]
  PIN eFPGA_result_b_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.056 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 47.5603 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 229.571 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 444.160000 550.160000 444.540000 ;
    END
  END eFPGA_result_b_i[1]
  PIN eFPGA_result_b_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5114 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.056 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 39.0048 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 179.849 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 447.820000 550.160000 448.200000 ;
    END
  END eFPGA_result_b_i[0]
  PIN eFPGA_result_c_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.784 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 50.0127 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 257.139 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 450.870000 550.160000 451.250000 ;
    END
  END eFPGA_result_c_i[31]
  PIN eFPGA_result_c_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.4498 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.536 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 25.9012 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 137.919 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 454.530000 550.160000 454.910000 ;
    END
  END eFPGA_result_c_i[30]
  PIN eFPGA_result_c_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.2948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 71.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 67.755 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 358.388 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 458.190000 550.160000 458.570000 ;
    END
  END eFPGA_result_c_i[29]
  PIN eFPGA_result_c_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.8438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.304 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 89.7634 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 471.188 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 461.240000 550.160000 461.620000 ;
    END
  END eFPGA_result_c_i[28]
  PIN eFPGA_result_c_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4846 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.816 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 25.2527 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 131.107 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 464.900000 550.160000 465.280000 ;
    END
  END eFPGA_result_c_i[27]
  PIN eFPGA_result_c_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.92 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 74.1618 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 369.313 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 468.560000 550.160000 468.940000 ;
    END
  END eFPGA_result_c_i[26]
  PIN eFPGA_result_c_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.0726 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 11.1194 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 61.3778 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 471.610000 550.160000 471.990000 ;
    END
  END eFPGA_result_c_i[25]
  PIN eFPGA_result_c_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.6938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.504 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 73.5226 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 375.895 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 475.270000 550.160000 475.650000 ;
    END
  END eFPGA_result_c_i[24]
  PIN eFPGA_result_c_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.488 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 71.1889 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 356.865 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 478.930000 550.160000 479.310000 ;
    END
  END eFPGA_result_c_i[23]
  PIN eFPGA_result_c_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0736 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.3078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 98.8091 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 518.444 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 481.980000 550.160000 482.360000 ;
    END
  END eFPGA_result_c_i[22]
  PIN eFPGA_result_c_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 12.7469 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 61.903 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 485.640000 550.160000 486.020000 ;
    END
  END eFPGA_result_c_i[21]
  PIN eFPGA_result_c_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.2546 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 87.632 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 83.5473 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 446.978 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 489.300000 550.160000 489.680000 ;
    END
  END eFPGA_result_c_i[20]
  PIN eFPGA_result_c_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 56.3897 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 279.931 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 492.350000 550.160000 492.730000 ;
    END
  END eFPGA_result_c_i[19]
  PIN eFPGA_result_c_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 13.9291 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 67.8141 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 496.010000 550.160000 496.390000 ;
    END
  END eFPGA_result_c_i[18]
  PIN eFPGA_result_c_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.864 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 13.256 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 65.1475 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 499.060000 550.160000 499.440000 ;
    END
  END eFPGA_result_c_i[17]
  PIN eFPGA_result_c_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.056 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 82.3008 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 413.737 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 502.720000 550.160000 503.100000 ;
    END
  END eFPGA_result_c_i[16]
  PIN eFPGA_result_c_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 77.6624 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 387.745 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 506.380000 550.160000 506.760000 ;
    END
  END eFPGA_result_c_i[15]
  PIN eFPGA_result_c_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 18.6547 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 91.2566 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 509.430000 550.160000 509.810000 ;
    END
  END eFPGA_result_c_i[14]
  PIN eFPGA_result_c_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 12.4616 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 60.1495 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 513.090000 550.160000 513.470000 ;
    END
  END eFPGA_result_c_i[13]
  PIN eFPGA_result_c_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 11.8572 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 56.8646 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 516.750000 550.160000 517.130000 ;
    END
  END eFPGA_result_c_i[12]
  PIN eFPGA_result_c_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.376 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 83.3877 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 419.345 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 519.800000 550.160000 520.180000 ;
    END
  END eFPGA_result_c_i[11]
  PIN eFPGA_result_c_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.442 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.96 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 12.2333 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 66.295 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 523.460000 550.160000 523.840000 ;
    END
  END eFPGA_result_c_i[10]
  PIN eFPGA_result_c_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 73.5978 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 365.774 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 527.120000 550.160000 527.500000 ;
    END
  END eFPGA_result_c_i[9]
  PIN eFPGA_result_c_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9624 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.128 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 7.28141 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 35.4465 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 530.170000 550.160000 530.550000 ;
    END
  END eFPGA_result_c_i[8]
  PIN eFPGA_result_c_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 14.9372 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 72.5939 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 533.830000 550.160000 534.210000 ;
    END
  END eFPGA_result_c_i[7]
  PIN eFPGA_result_c_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1674 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.888 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 61.163 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 307.697 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 537.490000 550.160000 537.870000 ;
    END
  END eFPGA_result_c_i[6]
  PIN eFPGA_result_c_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.704 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 83.016 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 416.307 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 540.540000 550.160000 540.920000 ;
    END
  END eFPGA_result_c_i[5]
  PIN eFPGA_result_c_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6524 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 23.5671 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 116.836 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 544.200000 550.160000 544.580000 ;
    END
  END eFPGA_result_c_i[4]
  PIN eFPGA_result_c_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6864 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.656 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 72.622 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 361.596 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 547.860000 550.160000 548.240000 ;
    END
  END eFPGA_result_c_i[3]
  PIN eFPGA_result_c_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7932 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.696 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 52.0543 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 265.046 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 550.910000 550.160000 551.290000 ;
    END
  END eFPGA_result_c_i[2]
  PIN eFPGA_result_c_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.28 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 77.4459 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 387.115 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 554.570000 550.160000 554.950000 ;
    END
  END eFPGA_result_c_i[1]
  PIN eFPGA_result_c_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.904 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 81.9897 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 411.984 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 558.230000 550.160000 558.610000 ;
    END
  END eFPGA_result_c_i[0]
  PIN eFPGA_write_strobe_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 561.280000 550.160000 561.660000 ;
    END
  END eFPGA_write_strobe_o
  PIN eFPGA_fpga_done_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.864 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 5.2901 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 26.0808 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 564.940000 550.160000 565.320000 ;
    END
  END eFPGA_fpga_done_i
  PIN eFPGA_en_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.5164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.416 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 568.600000 550.160000 568.980000 ;
    END
  END eFPGA_en_o
  PIN eFPGA_operator_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.448 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 571.650000 550.160000 572.030000 ;
    END
  END eFPGA_operator_o[1]
  PIN eFPGA_operator_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7726 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 58.4958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 312.448 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 575.310000 550.160000 575.690000 ;
    END
  END eFPGA_operator_o[0]
  PIN eFPGA_delay_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.4804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.224 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 578.970000 550.160000 579.350000 ;
    END
  END eFPGA_delay_o[3]
  PIN eFPGA_delay_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 582.020000 550.160000 582.400000 ;
    END
  END eFPGA_delay_o[2]
  PIN eFPGA_delay_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 585.680000 550.160000 586.060000 ;
    END
  END eFPGA_delay_o[1]
  PIN eFPGA_delay_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 549.260000 589.340000 550.160000 589.720000 ;
    END
  END eFPGA_delay_o[0]
  PIN irq_software_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0405 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.9198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 149.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 94.6364 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 501.479 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 345.040000 0.000000 345.420000 0.900000 ;
    END
  END irq_software_i
  PIN irq_timer_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8473 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.9826 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.848 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 11.9265 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 64.6748 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 346.420000 0.000000 346.800000 0.900000 ;
    END
  END irq_timer_i
  PIN irq_external_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7829 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.4066 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 157.776 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 77.7644 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 410.501 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 347.340000 0.000000 347.720000 0.900000 ;
    END
  END irq_external_i
  PIN irq_fast_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.113 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.339 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 6.47333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.1545 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 348.720000 0.000000 349.100000 0.900000 ;
    END
  END irq_fast_i[14]
  PIN irq_fast_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.253 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 10.1242 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 47.5182 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 350.100000 0.000000 350.480000 0.900000 ;
    END
  END irq_fast_i[13]
  PIN irq_fast_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1858 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.703 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.92909 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.4333 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 351.480000 0.000000 351.860000 0.900000 ;
    END
  END irq_fast_i[12]
  PIN irq_fast_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.666 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 6.83354 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 33.0919 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 352.860000 0.000000 353.240000 0.900000 ;
    END
  END irq_fast_i[11]
  PIN irq_fast_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6744 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.146 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 6.56667 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.6212 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 353.780000 0.000000 354.160000 0.900000 ;
    END
  END irq_fast_i[10]
  PIN irq_fast_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8808 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.168 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 8.77111 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 42.6232 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 355.160000 0.000000 355.540000 0.900000 ;
    END
  END irq_fast_i[9]
  PIN irq_fast_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.651 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.029 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 5.1497 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.5364 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 356.540000 0.000000 356.920000 0.900000 ;
    END
  END irq_fast_i[8]
  PIN irq_fast_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.1398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 129.216 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 58.0133 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 310.552 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 357.920000 0.000000 358.300000 0.900000 ;
    END
  END irq_fast_i[7]
  PIN irq_fast_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6121 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.8796 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 149.632 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 62.6865 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 334.475 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 358.840000 0.000000 359.220000 0.900000 ;
    END
  END irq_fast_i[6]
  PIN irq_fast_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3715 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.4605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.3916 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 109.696 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 49.1091 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 261.236 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 360.220000 0.000000 360.600000 0.900000 ;
    END
  END irq_fast_i[5]
  PIN irq_fast_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6058 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.803 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 5.67677 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 27.3081 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 361.600000 0.000000 361.980000 0.900000 ;
    END
  END irq_fast_i[4]
  PIN irq_fast_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8819 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.1305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.3286 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 93.36 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 48.1923 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 255.519 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 362.980000 0.000000 363.360000 0.900000 ;
    END
  END irq_fast_i[3]
  PIN irq_fast_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2499 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.9705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.9788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 91.024 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 55.3188 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 289.549 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 364.360000 0.000000 364.740000 0.900000 ;
    END
  END irq_fast_i[2]
  PIN irq_fast_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5629 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.717 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 5.86626 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 31.6909 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 365.280000 0.000000 365.660000 0.900000 ;
    END
  END irq_fast_i[1]
  PIN irq_fast_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.854 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.24395 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.0004 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 156.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 73.8319 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 396.079 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 366.660000 0.000000 367.040000 0.900000 ;
    END
  END irq_fast_i[0]
  PIN irq_nm_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8263 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.9705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.3442 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.384 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.873 LAYER met4  ;
    ANTENNAMAXAREACAR 53.7827 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 271.656 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32852 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 368.040000 0.000000 368.420000 0.900000 ;
    END
  END irq_nm_i
  PIN debug_req_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6917 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.18 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.76 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.3398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 105.968 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 65.2296 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 326.759 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.67778 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 369.420000 0.000000 369.800000 0.900000 ;
    END
  END debug_req_i
  PIN crash_dump_o[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.0516 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.914 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 370.800000 0.000000 371.180000 0.900000 ;
    END
  END crash_dump_o[127]
  PIN crash_dump_o[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4413 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.5668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 142.16 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 371.720000 0.000000 372.100000 0.900000 ;
    END
  END crash_dump_o[126]
  PIN crash_dump_o[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.0496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.022 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 373.100000 0.000000 373.480000 0.900000 ;
    END
  END crash_dump_o[125]
  PIN crash_dump_o[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0237 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.8395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.574 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.9158 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.688 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 374.480000 0.000000 374.860000 0.900000 ;
    END
  END crash_dump_o[124]
  PIN crash_dump_o[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9102 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.443 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 375.860000 0.000000 376.240000 0.900000 ;
    END
  END crash_dump_o[123]
  PIN crash_dump_o[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6034 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.791 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 376.780000 0.000000 377.160000 0.900000 ;
    END
  END crash_dump_o[122]
  PIN crash_dump_o[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.1946 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.747 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 378.160000 0.000000 378.540000 0.900000 ;
    END
  END crash_dump_o[121]
  PIN crash_dump_o[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6414 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.099 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 379.540000 0.000000 379.920000 0.900000 ;
    END
  END crash_dump_o[120]
  PIN crash_dump_o[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0264 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.863 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 38.0432 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 186.479 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via2  ;
    ANTENNADIFFAREA 4.5209 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.9828 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.712 LAYER met3  ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 54.1354 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 274.204 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 380.920000 0.000000 381.300000 0.900000 ;
    END
  END crash_dump_o[119]
  PIN crash_dump_o[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.4354 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.069 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 382.300000 0.000000 382.680000 0.900000 ;
    END
  END crash_dump_o[118]
  PIN crash_dump_o[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3722 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.753 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 383.220000 0.000000 383.600000 0.900000 ;
    END
  END crash_dump_o[117]
  PIN crash_dump_o[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.437 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 384.600000 0.000000 384.980000 0.900000 ;
    END
  END crash_dump_o[116]
  PIN crash_dump_o[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7142 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.345 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 385.980000 0.000000 386.360000 0.900000 ;
    END
  END crash_dump_o[115]
  PIN crash_dump_o[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.5402 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.475 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 387.360000 0.000000 387.740000 0.900000 ;
    END
  END crash_dump_o[114]
  PIN crash_dump_o[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1678 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.731 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 388.280000 0.000000 388.660000 0.900000 ;
    END
  END crash_dump_o[113]
  PIN crash_dump_o[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4064 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.914 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 389.660000 0.000000 390.040000 0.900000 ;
    END
  END crash_dump_o[112]
  PIN crash_dump_o[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.6266 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.025 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 391.040000 0.000000 391.420000 0.900000 ;
    END
  END crash_dump_o[111]
  PIN crash_dump_o[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4569 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.6938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.504 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 392.420000 0.000000 392.800000 0.900000 ;
    END
  END crash_dump_o[110]
  PIN crash_dump_o[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0218 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.001 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 393.800000 0.000000 394.180000 0.900000 ;
    END
  END crash_dump_o[109]
  PIN crash_dump_o[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.4998 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.391 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 394.720000 0.000000 395.100000 0.900000 ;
    END
  END crash_dump_o[108]
  PIN crash_dump_o[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.651 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.029 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 396.100000 0.000000 396.480000 0.900000 ;
    END
  END crash_dump_o[107]
  PIN crash_dump_o[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.0094 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.939 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 397.480000 0.000000 397.860000 0.900000 ;
    END
  END crash_dump_o[106]
  PIN crash_dump_o[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.949 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 398.860000 0.000000 399.240000 0.900000 ;
    END
  END crash_dump_o[105]
  PIN crash_dump_o[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.9758 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.771 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 399.780000 0.000000 400.160000 0.900000 ;
    END
  END crash_dump_o[104]
  PIN crash_dump_o[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.988 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 401.160000 0.000000 401.540000 0.900000 ;
    END
  END crash_dump_o[103]
  PIN crash_dump_o[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.6574 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.179 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 402.540000 0.000000 402.920000 0.900000 ;
    END
  END crash_dump_o[102]
  PIN crash_dump_o[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.277 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.277 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 403.920000 0.000000 404.300000 0.900000 ;
    END
  END crash_dump_o[101]
  PIN crash_dump_o[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.651 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.029 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 405.300000 0.000000 405.680000 0.900000 ;
    END
  END crash_dump_o[100]
  PIN crash_dump_o[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8418 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.983 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 406.220000 0.000000 406.600000 0.900000 ;
    END
  END crash_dump_o[99]
  PIN crash_dump_o[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9761 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.9088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 143.984 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 407.600000 0.000000 407.980000 0.900000 ;
    END
  END crash_dump_o[98]
  PIN crash_dump_o[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.9658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 96.288 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 408.980000 0.000000 409.360000 0.900000 ;
    END
  END crash_dump_o[97]
  PIN crash_dump_o[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9761 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.9024 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 134.224 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 410.360000 0.000000 410.740000 0.900000 ;
    END
  END crash_dump_o[96]
  PIN crash_dump_o[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.8978 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.381 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 411.280000 0.000000 411.660000 0.900000 ;
    END
  END crash_dump_o[95]
  PIN crash_dump_o[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3977 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.0638 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 86.144 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 412.660000 0.000000 413.040000 0.900000 ;
    END
  END crash_dump_o[94]
  PIN crash_dump_o[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.9568 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.558 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 414.040000 0.000000 414.420000 0.900000 ;
    END
  END crash_dump_o[93]
  PIN crash_dump_o[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5654 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.719 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 415.420000 0.000000 415.800000 0.900000 ;
    END
  END crash_dump_o[92]
  PIN crash_dump_o[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.0848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.256 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 416.800000 0.000000 417.180000 0.900000 ;
    END
  END crash_dump_o[91]
  PIN crash_dump_o[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.344 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 417.720000 0.000000 418.100000 0.900000 ;
    END
  END crash_dump_o[90]
  PIN crash_dump_o[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.9882 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.597 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 419.100000 0.000000 419.480000 0.900000 ;
    END
  END crash_dump_o[89]
  PIN crash_dump_o[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.4038 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 66.624 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 420.480000 0.000000 420.860000 0.900000 ;
    END
  END crash_dump_o[88]
  PIN crash_dump_o[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7789 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.125 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.4078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 141.312 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 421.860000 0.000000 422.240000 0.900000 ;
    END
  END crash_dump_o[87]
  PIN crash_dump_o[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.3196 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 141.312 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 423.240000 0.000000 423.620000 0.900000 ;
    END
  END crash_dump_o[86]
  PIN crash_dump_o[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.674 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.2948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 103.376 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 424.160000 0.000000 424.540000 0.900000 ;
    END
  END crash_dump_o[85]
  PIN crash_dump_o[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.678 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.3838 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 141.184 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 425.540000 0.000000 425.920000 0.900000 ;
    END
  END crash_dump_o[84]
  PIN crash_dump_o[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.039 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.087 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 426.920000 0.000000 427.300000 0.900000 ;
    END
  END crash_dump_o[83]
  PIN crash_dump_o[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6678 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.113 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 428.300000 0.000000 428.680000 0.900000 ;
    END
  END crash_dump_o[82]
  PIN crash_dump_o[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6678 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.113 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 429.220000 0.000000 429.600000 0.900000 ;
    END
  END crash_dump_o[81]
  PIN crash_dump_o[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8102 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 430.600000 0.000000 430.980000 0.900000 ;
    END
  END crash_dump_o[80]
  PIN crash_dump_o[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.4334 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.059 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 431.980000 0.000000 432.360000 0.900000 ;
    END
  END crash_dump_o[79]
  PIN crash_dump_o[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8006 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.895 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 433.360000 0.000000 433.740000 0.900000 ;
    END
  END crash_dump_o[78]
  PIN crash_dump_o[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3963 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.7484 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.736 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 434.740000 0.000000 435.120000 0.900000 ;
    END
  END crash_dump_o[77]
  PIN crash_dump_o[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.4718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.251 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 435.660000 0.000000 436.040000 0.900000 ;
    END
  END crash_dump_o[76]
  PIN crash_dump_o[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.669 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.119 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 437.040000 0.000000 437.420000 0.900000 ;
    END
  END crash_dump_o[75]
  PIN crash_dump_o[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.942 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.484 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 438.420000 0.000000 438.800000 0.900000 ;
    END
  END crash_dump_o[74]
  PIN crash_dump_o[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.9296 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 123.232 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 439.800000 0.000000 440.180000 0.900000 ;
    END
  END crash_dump_o[73]
  PIN crash_dump_o[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7016 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.282 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 440.720000 0.000000 441.100000 0.900000 ;
    END
  END crash_dump_o[72]
  PIN crash_dump_o[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.3502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.525 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 442.100000 0.000000 442.480000 0.900000 ;
    END
  END crash_dump_o[71]
  PIN crash_dump_o[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.359 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 443.480000 0.000000 443.860000 0.900000 ;
    END
  END crash_dump_o[70]
  PIN crash_dump_o[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.865 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.217 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 444.860000 0.000000 445.240000 0.900000 ;
    END
  END crash_dump_o[69]
  PIN crash_dump_o[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1982 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.883 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 446.240000 0.000000 446.620000 0.900000 ;
    END
  END crash_dump_o[68]
  PIN crash_dump_o[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6982 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.265 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 447.160000 0.000000 447.540000 0.900000 ;
    END
  END crash_dump_o[67]
  PIN crash_dump_o[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6989 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.006 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.0598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.456 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 448.540000 0.000000 448.920000 0.900000 ;
    END
  END crash_dump_o[66]
  PIN crash_dump_o[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.921 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 449.920000 0.000000 450.300000 0.900000 ;
    END
  END crash_dump_o[65]
  PIN crash_dump_o[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4629 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.9275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.597 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.984 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.284 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 121.2 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met4  ;
    ANTENNAMAXAREACAR 71.3594 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 367.233 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.622127 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 451.300000 0.000000 451.680000 0.900000 ;
    END
  END crash_dump_o[64]
  PIN crash_dump_o[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2533 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.1055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.7018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 142.88 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 452.220000 0.000000 452.600000 0.900000 ;
    END
  END crash_dump_o[63]
  PIN crash_dump_o[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3535 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.9328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 144.112 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 453.600000 0.000000 453.980000 0.900000 ;
    END
  END crash_dump_o[62]
  PIN crash_dump_o[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.5208 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 163.248 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 454.980000 0.000000 455.360000 0.900000 ;
    END
  END crash_dump_o[61]
  PIN crash_dump_o[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9151 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.86 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.4538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 88.224 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 456.360000 0.000000 456.740000 0.900000 ;
    END
  END crash_dump_o[60]
  PIN crash_dump_o[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3387 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.5325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.817 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.4558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 125.568 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 457.740000 0.000000 458.120000 0.900000 ;
    END
  END crash_dump_o[59]
  PIN crash_dump_o[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9349 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.746 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.8438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 106.304 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 458.660000 0.000000 459.040000 0.900000 ;
    END
  END crash_dump_o[58]
  PIN crash_dump_o[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9702 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.625 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 460.040000 0.000000 460.420000 0.900000 ;
    END
  END crash_dump_o[57]
  PIN crash_dump_o[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0143 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.972 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 106.984 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8568 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 101.04 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 461.420000 0.000000 461.800000 0.900000 ;
    END
  END crash_dump_o[56]
  PIN crash_dump_o[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0143 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.0048 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 112.496 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 462.800000 0.000000 463.180000 0.900000 ;
    END
  END crash_dump_o[55]
  PIN crash_dump_o[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.172 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.7096 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 127.392 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 463.720000 0.000000 464.100000 0.900000 ;
    END
  END crash_dump_o[54]
  PIN crash_dump_o[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4305 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.2378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 135.072 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 465.100000 0.000000 465.480000 0.900000 ;
    END
  END crash_dump_o[53]
  PIN crash_dump_o[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.3795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.747 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.9548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 90.896 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 466.480000 0.000000 466.860000 0.900000 ;
    END
  END crash_dump_o[52]
  PIN crash_dump_o[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6693 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.1855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.3578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 103.712 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 467.860000 0.000000 468.240000 0.900000 ;
    END
  END crash_dump_o[51]
  PIN crash_dump_o[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6445 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.0615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.6018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.68 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 469.240000 0.000000 469.620000 0.900000 ;
    END
  END crash_dump_o[50]
  PIN crash_dump_o[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7695 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.6865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.2508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 145.808 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 470.160000 0.000000 470.540000 0.900000 ;
    END
  END crash_dump_o[49]
  PIN crash_dump_o[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.781 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.4798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 109.696 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 471.540000 0.000000 471.920000 0.900000 ;
    END
  END crash_dump_o[48]
  PIN crash_dump_o[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2323 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.5286 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 163.76 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 472.920000 0.000000 473.300000 0.900000 ;
    END
  END crash_dump_o[47]
  PIN crash_dump_o[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8931 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.746 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.0748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.536 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 474.300000 0.000000 474.680000 0.900000 ;
    END
  END crash_dump_o[46]
  PIN crash_dump_o[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9403 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.5405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.278 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.2358 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 97.728 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 475.220000 0.000000 475.600000 0.900000 ;
    END
  END crash_dump_o[45]
  PIN crash_dump_o[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1431 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.229 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.1184 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 119.376 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 476.600000 0.000000 476.980000 0.900000 ;
    END
  END crash_dump_o[44]
  PIN crash_dump_o[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1755 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.7165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.231 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.3656 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 104.224 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 477.980000 0.000000 478.360000 0.900000 ;
    END
  END crash_dump_o[43]
  PIN crash_dump_o[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8931 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.1508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 102.608 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 479.360000 0.000000 479.740000 0.900000 ;
    END
  END crash_dump_o[42]
  PIN crash_dump_o[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1245 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.0686 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 214.64 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 480.740000 0.000000 481.120000 0.900000 ;
    END
  END crash_dump_o[41]
  PIN crash_dump_o[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4661 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.1695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.9906 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 150.224 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 481.660000 0.000000 482.040000 0.900000 ;
    END
  END crash_dump_o[40]
  PIN crash_dump_o[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8931 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.332 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.7368 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 116.4 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 483.040000 0.000000 483.420000 0.900000 ;
    END
  END crash_dump_o[39]
  PIN crash_dump_o[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7905 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.7915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.4646 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 280.752 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 484.420000 0.000000 484.800000 0.900000 ;
    END
  END crash_dump_o[38]
  PIN crash_dump_o[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4413 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.253 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.0406 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 155.824 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 485.800000 0.000000 486.180000 0.900000 ;
    END
  END crash_dump_o[37]
  PIN crash_dump_o[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.3155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.07 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.0308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 133.968 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 487.180000 0.000000 487.560000 0.900000 ;
    END
  END crash_dump_o[36]
  PIN crash_dump_o[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0143 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.16 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 66.6114 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 356.672 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 488.100000 0.000000 488.480000 0.900000 ;
    END
  END crash_dump_o[35]
  PIN crash_dump_o[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6803 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.3916 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 109.696 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 489.480000 0.000000 489.860000 0.900000 ;
    END
  END crash_dump_o[34]
  PIN crash_dump_o[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0143 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.4428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 98.832 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 490.860000 0.000000 491.240000 0.900000 ;
    END
  END crash_dump_o[33]
  PIN crash_dump_o[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6025 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.8515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.908 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.976 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.9878 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.072 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 492.240000 0.000000 492.620000 0.900000 ;
    END
  END crash_dump_o[32]
  PIN crash_dump_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1851 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.4338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 146.784 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 493.160000 0.000000 493.540000 0.900000 ;
    END
  END crash_dump_o[31]
  PIN crash_dump_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9575 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.6265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.6 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.7542 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 325.904 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 494.540000 0.000000 494.920000 0.900000 ;
    END
  END crash_dump_o[30]
  PIN crash_dump_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2347 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.0125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.783 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.976 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.0842 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 215.664 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 495.920000 0.000000 496.300000 0.900000 ;
    END
  END crash_dump_o[29]
  PIN crash_dump_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5515 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.5965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.4794 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 179.968 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 497.300000 0.000000 497.680000 0.900000 ;
    END
  END crash_dump_o[28]
  PIN crash_dump_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6975 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.0136 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 283.68 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 498.680000 0.000000 499.060000 0.900000 ;
    END
  END crash_dump_o[27]
  PIN crash_dump_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3387 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.5325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.47 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 87.9516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 470.016 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 499.600000 0.000000 499.980000 0.900000 ;
    END
  END crash_dump_o[26]
  PIN crash_dump_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9837 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.9268 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 64.08 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 500.980000 0.000000 501.360000 0.900000 ;
    END
  END crash_dump_o[25]
  PIN crash_dump_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.3225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.333 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.5566 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 206.576 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 502.360000 0.000000 502.740000 0.900000 ;
    END
  END crash_dump_o[24]
  PIN crash_dump_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8962 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.373 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 503.740000 0.000000 504.120000 0.900000 ;
    END
  END crash_dump_o[23]
  PIN crash_dump_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3917 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.6795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 79.2852 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 424.736 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 504.660000 0.000000 505.040000 0.900000 ;
    END
  END crash_dump_o[22]
  PIN crash_dump_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.332 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.0206 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 230.384 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 506.040000 0.000000 506.420000 0.900000 ;
    END
  END crash_dump_o[21]
  PIN crash_dump_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6582 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.183 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 507.420000 0.000000 507.800000 0.900000 ;
    END
  END crash_dump_o[20]
  PIN crash_dump_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0143 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 103.481 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 554.72 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 508.800000 0.000000 509.180000 0.900000 ;
    END
  END crash_dump_o[19]
  PIN crash_dump_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5895 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.242 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 200.976 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 510.180000 0.000000 510.560000 0.900000 ;
    END
  END crash_dump_o[18]
  PIN crash_dump_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1851 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.299 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 84.9738 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 456.016 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 511.100000 0.000000 511.480000 0.900000 ;
    END
  END crash_dump_o[17]
  PIN crash_dump_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 120.946 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 646.928 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 512.480000 0.000000 512.860000 0.900000 ;
    END
  END crash_dump_o[16]
  PIN crash_dump_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 178.169 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 953.056 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 513.860000 0.000000 514.240000 0.900000 ;
    END
  END crash_dump_o[15]
  PIN crash_dump_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1431 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 145.151 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 775.552 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 515.240000 0.000000 515.620000 0.900000 ;
    END
  END crash_dump_o[14]
  PIN crash_dump_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0219 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.9485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 166.617 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 890.976 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 516.160000 0.000000 516.540000 0.900000 ;
    END
  END crash_dump_o[13]
  PIN crash_dump_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6159 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.9185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.782 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 159.233 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 852.064 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 517.540000 0.000000 517.920000 0.900000 ;
    END
  END crash_dump_o[12]
  PIN crash_dump_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2785 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.1135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.436 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 67.581 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 362.784 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 518.920000 0.000000 519.300000 0.900000 ;
    END
  END crash_dump_o[11]
  PIN crash_dump_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1245 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 108.112 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 578.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 520.300000 0.000000 520.680000 0.900000 ;
    END
  END crash_dump_o[10]
  PIN crash_dump_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9746 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.765 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 521.680000 0.000000 522.060000 0.900000 ;
    END
  END crash_dump_o[9]
  PIN crash_dump_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6582 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.183 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 522.600000 0.000000 522.980000 0.900000 ;
    END
  END crash_dump_o[8]
  PIN crash_dump_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.7764 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 327.904 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 523.980000 0.000000 524.360000 0.900000 ;
    END
  END crash_dump_o[7]
  PIN crash_dump_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 100.314 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 537.36 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 525.360000 0.000000 525.740000 0.900000 ;
    END
  END crash_dump_o[6]
  PIN crash_dump_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7905 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.7915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 102.717 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 550.176 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 526.740000 0.000000 527.120000 0.900000 ;
    END
  END crash_dump_o[5]
  PIN crash_dump_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.1035 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.3465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.046 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 71.559 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 384 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 527.660000 0.000000 528.040000 0.900000 ;
    END
  END crash_dump_o[4]
  PIN crash_dump_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 103.919 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 555.648 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 529.040000 0.000000 529.420000 0.900000 ;
    END
  END crash_dump_o[3]
  PIN crash_dump_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6443 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.9425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.3758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.808 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 530.420000 0.000000 530.800000 0.900000 ;
    END
  END crash_dump_o[2]
  PIN crash_dump_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0997 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.299 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 170.873 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 914.144 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 531.800000 0.000000 532.180000 0.900000 ;
    END
  END crash_dump_o[1]
  PIN crash_dump_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.2007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.8425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.84 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.8102 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 107.536 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 533.180000 0.000000 533.560000 0.900000 ;
    END
  END crash_dump_o[0]
  PIN fetch_enable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 37.0768 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 201.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.8542 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.104 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 57.6024 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 311.738 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 534.100000 0.000000 534.480000 0.900000 ;
    END
  END fetch_enable_i
  PIN alert_minor_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9578 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.681 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 535.480000 0.000000 535.860000 0.900000 ;
    END
  END alert_minor_o
  PIN alert_major_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8088 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.784 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 536.860000 0.000000 537.240000 0.900000 ;
    END
  END alert_major_o
  PIN core_sleep_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.906 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.52 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 538.240000 0.000000 538.620000 0.900000 ;
    END
  END core_sleep_o
  PIN scan_rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.160000 0.000000 539.540000 0.900000 ;
    END
  END scan_rst_ni
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 548.960000 592.790000 550.160000 593.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 592.790000 1.200000 593.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 548.960000 5.430000 550.160000 6.630000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 5.430000 1.200000 6.630000 ;
    END
    PORT
      LAYER met4 ;
        RECT 543.400000 598.560000 544.600000 599.760000 ;
    END
    PORT
      LAYER met4 ;
        RECT 543.400000 0.000000 544.600000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 5.560000 598.560000 6.760000 599.760000 ;
    END
    PORT
      LAYER met4 ;
        RECT 5.560000 0.000000 6.760000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 5.430000 550.160000 6.630000 ;
        RECT 0.000000 592.790000 550.160000 593.990000 ;
        RECT 5.560000 74.900000 6.760000 75.380000 ;
        RECT 102.120000 74.900000 103.320000 75.380000 ;
        RECT 57.120000 74.900000 58.320000 75.380000 ;
        RECT 12.120000 74.900000 13.320000 75.380000 ;
        RECT 12.120000 9.620000 13.320000 10.100000 ;
        RECT 12.120000 15.060000 13.320000 15.540000 ;
        RECT 12.120000 20.500000 13.320000 20.980000 ;
        RECT 12.120000 25.940000 13.320000 26.420000 ;
        RECT 12.120000 31.380000 13.320000 31.860000 ;
        RECT 12.120000 36.820000 13.320000 37.300000 ;
        RECT 5.560000 9.620000 6.760000 10.100000 ;
        RECT 5.560000 15.060000 6.760000 15.540000 ;
        RECT 5.560000 20.500000 6.760000 20.980000 ;
        RECT 5.560000 25.940000 6.760000 26.420000 ;
        RECT 5.560000 36.820000 6.760000 37.300000 ;
        RECT 5.560000 31.380000 6.760000 31.860000 ;
        RECT 12.120000 69.460000 13.320000 69.940000 ;
        RECT 12.120000 64.020000 13.320000 64.500000 ;
        RECT 12.120000 58.580000 13.320000 59.060000 ;
        RECT 12.120000 42.260000 13.320000 42.740000 ;
        RECT 12.120000 47.700000 13.320000 48.180000 ;
        RECT 12.120000 53.140000 13.320000 53.620000 ;
        RECT 5.560000 42.260000 6.760000 42.740000 ;
        RECT 5.560000 47.700000 6.760000 48.180000 ;
        RECT 5.560000 53.140000 6.760000 53.620000 ;
        RECT 5.560000 58.580000 6.760000 59.060000 ;
        RECT 5.560000 64.020000 6.760000 64.500000 ;
        RECT 5.560000 69.460000 6.760000 69.940000 ;
        RECT 57.120000 9.620000 58.320000 10.100000 ;
        RECT 57.120000 15.060000 58.320000 15.540000 ;
        RECT 57.120000 20.500000 58.320000 20.980000 ;
        RECT 57.120000 25.940000 58.320000 26.420000 ;
        RECT 57.120000 31.380000 58.320000 31.860000 ;
        RECT 57.120000 36.820000 58.320000 37.300000 ;
        RECT 102.120000 9.620000 103.320000 10.100000 ;
        RECT 102.120000 15.060000 103.320000 15.540000 ;
        RECT 102.120000 20.500000 103.320000 20.980000 ;
        RECT 102.120000 25.940000 103.320000 26.420000 ;
        RECT 102.120000 31.380000 103.320000 31.860000 ;
        RECT 102.120000 36.820000 103.320000 37.300000 ;
        RECT 57.120000 53.140000 58.320000 53.620000 ;
        RECT 57.120000 47.700000 58.320000 48.180000 ;
        RECT 57.120000 42.260000 58.320000 42.740000 ;
        RECT 57.120000 64.020000 58.320000 64.500000 ;
        RECT 57.120000 58.580000 58.320000 59.060000 ;
        RECT 57.120000 69.460000 58.320000 69.940000 ;
        RECT 102.120000 53.140000 103.320000 53.620000 ;
        RECT 102.120000 47.700000 103.320000 48.180000 ;
        RECT 102.120000 42.260000 103.320000 42.740000 ;
        RECT 102.120000 64.020000 103.320000 64.500000 ;
        RECT 102.120000 58.580000 103.320000 59.060000 ;
        RECT 102.120000 69.460000 103.320000 69.940000 ;
        RECT 12.120000 96.660000 13.320000 97.140000 ;
        RECT 12.120000 91.220000 13.320000 91.700000 ;
        RECT 12.120000 85.780000 13.320000 86.260000 ;
        RECT 12.120000 80.340000 13.320000 80.820000 ;
        RECT 12.120000 102.100000 13.320000 102.580000 ;
        RECT 12.120000 107.540000 13.320000 108.020000 ;
        RECT 5.560000 80.340000 6.760000 80.820000 ;
        RECT 5.560000 85.780000 6.760000 86.260000 ;
        RECT 5.560000 91.220000 6.760000 91.700000 ;
        RECT 5.560000 96.660000 6.760000 97.140000 ;
        RECT 5.560000 102.100000 6.760000 102.580000 ;
        RECT 5.560000 107.540000 6.760000 108.020000 ;
        RECT 12.120000 145.620000 13.320000 146.100000 ;
        RECT 12.120000 140.180000 13.320000 140.660000 ;
        RECT 12.120000 134.740000 13.320000 135.220000 ;
        RECT 12.120000 112.980000 13.320000 113.460000 ;
        RECT 12.120000 118.420000 13.320000 118.900000 ;
        RECT 12.120000 123.860000 13.320000 124.340000 ;
        RECT 12.120000 129.300000 13.320000 129.780000 ;
        RECT 5.560000 112.980000 6.760000 113.460000 ;
        RECT 5.560000 118.420000 6.760000 118.900000 ;
        RECT 5.560000 123.860000 6.760000 124.340000 ;
        RECT 5.560000 129.300000 6.760000 129.780000 ;
        RECT 5.560000 140.180000 6.760000 140.660000 ;
        RECT 5.560000 134.740000 6.760000 135.220000 ;
        RECT 5.560000 145.620000 6.760000 146.100000 ;
        RECT 57.120000 91.220000 58.320000 91.700000 ;
        RECT 57.120000 85.780000 58.320000 86.260000 ;
        RECT 57.120000 80.340000 58.320000 80.820000 ;
        RECT 57.120000 107.540000 58.320000 108.020000 ;
        RECT 57.120000 96.660000 58.320000 97.140000 ;
        RECT 57.120000 102.100000 58.320000 102.580000 ;
        RECT 102.120000 91.220000 103.320000 91.700000 ;
        RECT 102.120000 85.780000 103.320000 86.260000 ;
        RECT 102.120000 80.340000 103.320000 80.820000 ;
        RECT 102.120000 96.660000 103.320000 97.140000 ;
        RECT 102.120000 102.100000 103.320000 102.580000 ;
        RECT 102.120000 107.540000 103.320000 108.020000 ;
        RECT 57.120000 129.300000 58.320000 129.780000 ;
        RECT 57.120000 123.860000 58.320000 124.340000 ;
        RECT 57.120000 118.420000 58.320000 118.900000 ;
        RECT 57.120000 112.980000 58.320000 113.460000 ;
        RECT 57.120000 134.740000 58.320000 135.220000 ;
        RECT 57.120000 140.180000 58.320000 140.660000 ;
        RECT 57.120000 145.620000 58.320000 146.100000 ;
        RECT 102.120000 129.300000 103.320000 129.780000 ;
        RECT 102.120000 123.860000 103.320000 124.340000 ;
        RECT 102.120000 118.420000 103.320000 118.900000 ;
        RECT 102.120000 112.980000 103.320000 113.460000 ;
        RECT 102.120000 134.740000 103.320000 135.220000 ;
        RECT 102.120000 140.180000 103.320000 140.660000 ;
        RECT 102.120000 145.620000 103.320000 146.100000 ;
        RECT 192.120000 74.900000 193.320000 75.380000 ;
        RECT 147.120000 74.900000 148.320000 75.380000 ;
        RECT 237.120000 74.900000 238.320000 75.380000 ;
        RECT 147.120000 9.620000 148.320000 10.100000 ;
        RECT 147.120000 15.060000 148.320000 15.540000 ;
        RECT 147.120000 20.500000 148.320000 20.980000 ;
        RECT 147.120000 25.940000 148.320000 26.420000 ;
        RECT 147.120000 31.380000 148.320000 31.860000 ;
        RECT 147.120000 36.820000 148.320000 37.300000 ;
        RECT 192.120000 9.620000 193.320000 10.100000 ;
        RECT 192.120000 15.060000 193.320000 15.540000 ;
        RECT 192.120000 20.500000 193.320000 20.980000 ;
        RECT 192.120000 25.940000 193.320000 26.420000 ;
        RECT 192.120000 31.380000 193.320000 31.860000 ;
        RECT 192.120000 36.820000 193.320000 37.300000 ;
        RECT 147.120000 53.140000 148.320000 53.620000 ;
        RECT 147.120000 47.700000 148.320000 48.180000 ;
        RECT 147.120000 42.260000 148.320000 42.740000 ;
        RECT 147.120000 64.020000 148.320000 64.500000 ;
        RECT 147.120000 58.580000 148.320000 59.060000 ;
        RECT 147.120000 69.460000 148.320000 69.940000 ;
        RECT 192.120000 53.140000 193.320000 53.620000 ;
        RECT 192.120000 47.700000 193.320000 48.180000 ;
        RECT 192.120000 42.260000 193.320000 42.740000 ;
        RECT 192.120000 64.020000 193.320000 64.500000 ;
        RECT 192.120000 58.580000 193.320000 59.060000 ;
        RECT 192.120000 69.460000 193.320000 69.940000 ;
        RECT 237.120000 9.620000 238.320000 10.100000 ;
        RECT 237.120000 15.060000 238.320000 15.540000 ;
        RECT 237.120000 20.500000 238.320000 20.980000 ;
        RECT 237.120000 25.940000 238.320000 26.420000 ;
        RECT 237.120000 31.380000 238.320000 31.860000 ;
        RECT 237.120000 36.820000 238.320000 37.300000 ;
        RECT 237.120000 69.460000 238.320000 69.940000 ;
        RECT 237.120000 64.020000 238.320000 64.500000 ;
        RECT 237.120000 42.260000 238.320000 42.740000 ;
        RECT 237.120000 47.700000 238.320000 48.180000 ;
        RECT 237.120000 53.140000 238.320000 53.620000 ;
        RECT 237.120000 58.580000 238.320000 59.060000 ;
        RECT 147.120000 91.220000 148.320000 91.700000 ;
        RECT 147.120000 85.780000 148.320000 86.260000 ;
        RECT 147.120000 80.340000 148.320000 80.820000 ;
        RECT 147.120000 107.540000 148.320000 108.020000 ;
        RECT 147.120000 96.660000 148.320000 97.140000 ;
        RECT 147.120000 102.100000 148.320000 102.580000 ;
        RECT 192.120000 91.220000 193.320000 91.700000 ;
        RECT 192.120000 85.780000 193.320000 86.260000 ;
        RECT 192.120000 80.340000 193.320000 80.820000 ;
        RECT 192.120000 96.660000 193.320000 97.140000 ;
        RECT 192.120000 102.100000 193.320000 102.580000 ;
        RECT 192.120000 107.540000 193.320000 108.020000 ;
        RECT 147.120000 129.300000 148.320000 129.780000 ;
        RECT 147.120000 123.860000 148.320000 124.340000 ;
        RECT 147.120000 118.420000 148.320000 118.900000 ;
        RECT 147.120000 112.980000 148.320000 113.460000 ;
        RECT 147.120000 134.740000 148.320000 135.220000 ;
        RECT 147.120000 140.180000 148.320000 140.660000 ;
        RECT 147.120000 145.620000 148.320000 146.100000 ;
        RECT 192.120000 129.300000 193.320000 129.780000 ;
        RECT 192.120000 123.860000 193.320000 124.340000 ;
        RECT 192.120000 118.420000 193.320000 118.900000 ;
        RECT 192.120000 112.980000 193.320000 113.460000 ;
        RECT 192.120000 134.740000 193.320000 135.220000 ;
        RECT 192.120000 140.180000 193.320000 140.660000 ;
        RECT 192.120000 145.620000 193.320000 146.100000 ;
        RECT 237.120000 96.660000 238.320000 97.140000 ;
        RECT 237.120000 91.220000 238.320000 91.700000 ;
        RECT 237.120000 85.780000 238.320000 86.260000 ;
        RECT 237.120000 80.340000 238.320000 80.820000 ;
        RECT 237.120000 102.100000 238.320000 102.580000 ;
        RECT 237.120000 107.540000 238.320000 108.020000 ;
        RECT 237.120000 145.620000 238.320000 146.100000 ;
        RECT 237.120000 140.180000 238.320000 140.660000 ;
        RECT 237.120000 134.740000 238.320000 135.220000 ;
        RECT 237.120000 112.980000 238.320000 113.460000 ;
        RECT 237.120000 118.420000 238.320000 118.900000 ;
        RECT 237.120000 123.860000 238.320000 124.340000 ;
        RECT 237.120000 129.300000 238.320000 129.780000 ;
        RECT 12.120000 156.500000 13.320000 156.980000 ;
        RECT 12.120000 151.060000 13.320000 151.540000 ;
        RECT 12.120000 161.940000 13.320000 162.420000 ;
        RECT 12.120000 167.380000 13.320000 167.860000 ;
        RECT 12.120000 172.820000 13.320000 173.300000 ;
        RECT 12.120000 178.260000 13.320000 178.740000 ;
        RECT 12.120000 183.700000 13.320000 184.180000 ;
        RECT 5.560000 151.060000 6.760000 151.540000 ;
        RECT 5.560000 156.500000 6.760000 156.980000 ;
        RECT 5.560000 161.940000 6.760000 162.420000 ;
        RECT 5.560000 167.380000 6.760000 167.860000 ;
        RECT 5.560000 172.820000 6.760000 173.300000 ;
        RECT 5.560000 183.700000 6.760000 184.180000 ;
        RECT 5.560000 178.260000 6.760000 178.740000 ;
        RECT 12.120000 221.780000 13.320000 222.260000 ;
        RECT 12.120000 216.340000 13.320000 216.820000 ;
        RECT 12.120000 210.900000 13.320000 211.380000 ;
        RECT 12.120000 205.460000 13.320000 205.940000 ;
        RECT 12.120000 189.140000 13.320000 189.620000 ;
        RECT 12.120000 194.580000 13.320000 195.060000 ;
        RECT 12.120000 200.020000 13.320000 200.500000 ;
        RECT 5.560000 189.140000 6.760000 189.620000 ;
        RECT 5.560000 194.580000 6.760000 195.060000 ;
        RECT 5.560000 200.020000 6.760000 200.500000 ;
        RECT 5.560000 205.460000 6.760000 205.940000 ;
        RECT 5.560000 210.900000 6.760000 211.380000 ;
        RECT 5.560000 221.780000 6.760000 222.260000 ;
        RECT 5.560000 216.340000 6.760000 216.820000 ;
        RECT 57.120000 167.380000 58.320000 167.860000 ;
        RECT 57.120000 156.500000 58.320000 156.980000 ;
        RECT 57.120000 151.060000 58.320000 151.540000 ;
        RECT 57.120000 161.940000 58.320000 162.420000 ;
        RECT 57.120000 178.260000 58.320000 178.740000 ;
        RECT 57.120000 172.820000 58.320000 173.300000 ;
        RECT 57.120000 183.700000 58.320000 184.180000 ;
        RECT 102.120000 156.500000 103.320000 156.980000 ;
        RECT 102.120000 151.060000 103.320000 151.540000 ;
        RECT 102.120000 161.940000 103.320000 162.420000 ;
        RECT 102.120000 167.380000 103.320000 167.860000 ;
        RECT 102.120000 172.820000 103.320000 173.300000 ;
        RECT 102.120000 178.260000 103.320000 178.740000 ;
        RECT 102.120000 183.700000 103.320000 184.180000 ;
        RECT 57.120000 205.460000 58.320000 205.940000 ;
        RECT 57.120000 200.020000 58.320000 200.500000 ;
        RECT 57.120000 194.580000 58.320000 195.060000 ;
        RECT 57.120000 189.140000 58.320000 189.620000 ;
        RECT 57.120000 210.900000 58.320000 211.380000 ;
        RECT 57.120000 216.340000 58.320000 216.820000 ;
        RECT 57.120000 221.780000 58.320000 222.260000 ;
        RECT 102.120000 205.460000 103.320000 205.940000 ;
        RECT 102.120000 200.020000 103.320000 200.500000 ;
        RECT 102.120000 194.580000 103.320000 195.060000 ;
        RECT 102.120000 189.140000 103.320000 189.620000 ;
        RECT 102.120000 210.900000 103.320000 211.380000 ;
        RECT 102.120000 216.340000 103.320000 216.820000 ;
        RECT 102.120000 221.780000 103.320000 222.260000 ;
        RECT 12.120000 243.540000 13.320000 244.020000 ;
        RECT 12.120000 238.100000 13.320000 238.580000 ;
        RECT 12.120000 232.660000 13.320000 233.140000 ;
        RECT 12.120000 227.220000 13.320000 227.700000 ;
        RECT 12.120000 248.980000 13.320000 249.460000 ;
        RECT 12.120000 254.420000 13.320000 254.900000 ;
        RECT 12.120000 259.860000 13.320000 260.340000 ;
        RECT 5.560000 243.540000 6.760000 244.020000 ;
        RECT 5.560000 227.220000 6.760000 227.700000 ;
        RECT 5.560000 232.660000 6.760000 233.140000 ;
        RECT 5.560000 238.100000 6.760000 238.580000 ;
        RECT 5.560000 248.980000 6.760000 249.460000 ;
        RECT 5.560000 259.860000 6.760000 260.340000 ;
        RECT 5.560000 254.420000 6.760000 254.900000 ;
        RECT 12.120000 297.940000 13.320000 298.420000 ;
        RECT 12.120000 292.500000 13.320000 292.980000 ;
        RECT 12.120000 287.060000 13.320000 287.540000 ;
        RECT 12.120000 281.620000 13.320000 282.100000 ;
        RECT 12.120000 265.300000 13.320000 265.780000 ;
        RECT 12.120000 270.740000 13.320000 271.220000 ;
        RECT 12.120000 276.180000 13.320000 276.660000 ;
        RECT 5.560000 265.300000 6.760000 265.780000 ;
        RECT 5.560000 270.740000 6.760000 271.220000 ;
        RECT 5.560000 276.180000 6.760000 276.660000 ;
        RECT 5.560000 281.620000 6.760000 282.100000 ;
        RECT 5.560000 287.060000 6.760000 287.540000 ;
        RECT 5.560000 297.940000 6.760000 298.420000 ;
        RECT 5.560000 292.500000 6.760000 292.980000 ;
        RECT 57.120000 243.540000 58.320000 244.020000 ;
        RECT 57.120000 238.100000 58.320000 238.580000 ;
        RECT 57.120000 232.660000 58.320000 233.140000 ;
        RECT 57.120000 227.220000 58.320000 227.700000 ;
        RECT 57.120000 254.420000 58.320000 254.900000 ;
        RECT 57.120000 248.980000 58.320000 249.460000 ;
        RECT 57.120000 259.860000 58.320000 260.340000 ;
        RECT 102.120000 243.540000 103.320000 244.020000 ;
        RECT 102.120000 238.100000 103.320000 238.580000 ;
        RECT 102.120000 232.660000 103.320000 233.140000 ;
        RECT 102.120000 227.220000 103.320000 227.700000 ;
        RECT 102.120000 248.980000 103.320000 249.460000 ;
        RECT 102.120000 254.420000 103.320000 254.900000 ;
        RECT 102.120000 259.860000 103.320000 260.340000 ;
        RECT 57.120000 276.180000 58.320000 276.660000 ;
        RECT 57.120000 270.740000 58.320000 271.220000 ;
        RECT 57.120000 265.300000 58.320000 265.780000 ;
        RECT 57.120000 287.060000 58.320000 287.540000 ;
        RECT 57.120000 281.620000 58.320000 282.100000 ;
        RECT 57.120000 292.500000 58.320000 292.980000 ;
        RECT 57.120000 297.940000 58.320000 298.420000 ;
        RECT 102.120000 276.180000 103.320000 276.660000 ;
        RECT 102.120000 270.740000 103.320000 271.220000 ;
        RECT 102.120000 265.300000 103.320000 265.780000 ;
        RECT 102.120000 287.060000 103.320000 287.540000 ;
        RECT 102.120000 281.620000 103.320000 282.100000 ;
        RECT 102.120000 292.500000 103.320000 292.980000 ;
        RECT 102.120000 297.940000 103.320000 298.420000 ;
        RECT 147.120000 167.380000 148.320000 167.860000 ;
        RECT 147.120000 151.060000 148.320000 151.540000 ;
        RECT 147.120000 156.500000 148.320000 156.980000 ;
        RECT 147.120000 161.940000 148.320000 162.420000 ;
        RECT 147.120000 178.260000 148.320000 178.740000 ;
        RECT 147.120000 172.820000 148.320000 173.300000 ;
        RECT 147.120000 183.700000 148.320000 184.180000 ;
        RECT 192.120000 151.060000 193.320000 151.540000 ;
        RECT 192.120000 156.500000 193.320000 156.980000 ;
        RECT 192.120000 161.940000 193.320000 162.420000 ;
        RECT 192.120000 167.380000 193.320000 167.860000 ;
        RECT 192.120000 172.820000 193.320000 173.300000 ;
        RECT 192.120000 178.260000 193.320000 178.740000 ;
        RECT 192.120000 183.700000 193.320000 184.180000 ;
        RECT 147.120000 205.460000 148.320000 205.940000 ;
        RECT 147.120000 200.020000 148.320000 200.500000 ;
        RECT 147.120000 194.580000 148.320000 195.060000 ;
        RECT 147.120000 189.140000 148.320000 189.620000 ;
        RECT 147.120000 210.900000 148.320000 211.380000 ;
        RECT 147.120000 216.340000 148.320000 216.820000 ;
        RECT 147.120000 221.780000 148.320000 222.260000 ;
        RECT 192.120000 205.460000 193.320000 205.940000 ;
        RECT 192.120000 200.020000 193.320000 200.500000 ;
        RECT 192.120000 194.580000 193.320000 195.060000 ;
        RECT 192.120000 189.140000 193.320000 189.620000 ;
        RECT 192.120000 210.900000 193.320000 211.380000 ;
        RECT 192.120000 216.340000 193.320000 216.820000 ;
        RECT 192.120000 221.780000 193.320000 222.260000 ;
        RECT 237.120000 156.500000 238.320000 156.980000 ;
        RECT 237.120000 151.060000 238.320000 151.540000 ;
        RECT 237.120000 161.940000 238.320000 162.420000 ;
        RECT 237.120000 167.380000 238.320000 167.860000 ;
        RECT 237.120000 172.820000 238.320000 173.300000 ;
        RECT 237.120000 178.260000 238.320000 178.740000 ;
        RECT 237.120000 183.700000 238.320000 184.180000 ;
        RECT 237.120000 221.780000 238.320000 222.260000 ;
        RECT 237.120000 216.340000 238.320000 216.820000 ;
        RECT 237.120000 210.900000 238.320000 211.380000 ;
        RECT 237.120000 205.460000 238.320000 205.940000 ;
        RECT 237.120000 189.140000 238.320000 189.620000 ;
        RECT 237.120000 194.580000 238.320000 195.060000 ;
        RECT 237.120000 200.020000 238.320000 200.500000 ;
        RECT 147.120000 243.540000 148.320000 244.020000 ;
        RECT 147.120000 238.100000 148.320000 238.580000 ;
        RECT 147.120000 232.660000 148.320000 233.140000 ;
        RECT 147.120000 227.220000 148.320000 227.700000 ;
        RECT 147.120000 254.420000 148.320000 254.900000 ;
        RECT 147.120000 248.980000 148.320000 249.460000 ;
        RECT 147.120000 259.860000 148.320000 260.340000 ;
        RECT 192.120000 243.540000 193.320000 244.020000 ;
        RECT 192.120000 238.100000 193.320000 238.580000 ;
        RECT 192.120000 232.660000 193.320000 233.140000 ;
        RECT 192.120000 227.220000 193.320000 227.700000 ;
        RECT 192.120000 248.980000 193.320000 249.460000 ;
        RECT 192.120000 254.420000 193.320000 254.900000 ;
        RECT 192.120000 259.860000 193.320000 260.340000 ;
        RECT 147.120000 276.180000 148.320000 276.660000 ;
        RECT 147.120000 270.740000 148.320000 271.220000 ;
        RECT 147.120000 265.300000 148.320000 265.780000 ;
        RECT 147.120000 287.060000 148.320000 287.540000 ;
        RECT 147.120000 281.620000 148.320000 282.100000 ;
        RECT 147.120000 292.500000 148.320000 292.980000 ;
        RECT 147.120000 297.940000 148.320000 298.420000 ;
        RECT 192.120000 276.180000 193.320000 276.660000 ;
        RECT 192.120000 270.740000 193.320000 271.220000 ;
        RECT 192.120000 265.300000 193.320000 265.780000 ;
        RECT 192.120000 287.060000 193.320000 287.540000 ;
        RECT 192.120000 281.620000 193.320000 282.100000 ;
        RECT 192.120000 292.500000 193.320000 292.980000 ;
        RECT 192.120000 297.940000 193.320000 298.420000 ;
        RECT 237.120000 243.540000 238.320000 244.020000 ;
        RECT 237.120000 238.100000 238.320000 238.580000 ;
        RECT 237.120000 232.660000 238.320000 233.140000 ;
        RECT 237.120000 227.220000 238.320000 227.700000 ;
        RECT 237.120000 248.980000 238.320000 249.460000 ;
        RECT 237.120000 254.420000 238.320000 254.900000 ;
        RECT 237.120000 259.860000 238.320000 260.340000 ;
        RECT 237.120000 297.940000 238.320000 298.420000 ;
        RECT 237.120000 292.500000 238.320000 292.980000 ;
        RECT 237.120000 287.060000 238.320000 287.540000 ;
        RECT 237.120000 281.620000 238.320000 282.100000 ;
        RECT 237.120000 265.300000 238.320000 265.780000 ;
        RECT 237.120000 270.740000 238.320000 271.220000 ;
        RECT 237.120000 276.180000 238.320000 276.660000 ;
        RECT 417.120000 74.900000 418.320000 75.380000 ;
        RECT 372.120000 74.900000 373.320000 75.380000 ;
        RECT 327.120000 74.900000 328.320000 75.380000 ;
        RECT 282.120000 74.900000 283.320000 75.380000 ;
        RECT 282.120000 9.620000 283.320000 10.100000 ;
        RECT 282.120000 15.060000 283.320000 15.540000 ;
        RECT 282.120000 20.500000 283.320000 20.980000 ;
        RECT 282.120000 25.940000 283.320000 26.420000 ;
        RECT 282.120000 31.380000 283.320000 31.860000 ;
        RECT 282.120000 36.820000 283.320000 37.300000 ;
        RECT 327.120000 9.620000 328.320000 10.100000 ;
        RECT 327.120000 15.060000 328.320000 15.540000 ;
        RECT 327.120000 20.500000 328.320000 20.980000 ;
        RECT 327.120000 25.940000 328.320000 26.420000 ;
        RECT 327.120000 31.380000 328.320000 31.860000 ;
        RECT 327.120000 36.820000 328.320000 37.300000 ;
        RECT 282.120000 53.140000 283.320000 53.620000 ;
        RECT 282.120000 47.700000 283.320000 48.180000 ;
        RECT 282.120000 42.260000 283.320000 42.740000 ;
        RECT 282.120000 64.020000 283.320000 64.500000 ;
        RECT 282.120000 58.580000 283.320000 59.060000 ;
        RECT 282.120000 69.460000 283.320000 69.940000 ;
        RECT 327.120000 53.140000 328.320000 53.620000 ;
        RECT 327.120000 47.700000 328.320000 48.180000 ;
        RECT 327.120000 42.260000 328.320000 42.740000 ;
        RECT 327.120000 64.020000 328.320000 64.500000 ;
        RECT 327.120000 58.580000 328.320000 59.060000 ;
        RECT 327.120000 69.460000 328.320000 69.940000 ;
        RECT 372.120000 9.620000 373.320000 10.100000 ;
        RECT 372.120000 15.060000 373.320000 15.540000 ;
        RECT 372.120000 20.500000 373.320000 20.980000 ;
        RECT 372.120000 25.940000 373.320000 26.420000 ;
        RECT 372.120000 31.380000 373.320000 31.860000 ;
        RECT 372.120000 36.820000 373.320000 37.300000 ;
        RECT 417.120000 9.620000 418.320000 10.100000 ;
        RECT 417.120000 15.060000 418.320000 15.540000 ;
        RECT 417.120000 20.500000 418.320000 20.980000 ;
        RECT 417.120000 25.940000 418.320000 26.420000 ;
        RECT 417.120000 31.380000 418.320000 31.860000 ;
        RECT 417.120000 36.820000 418.320000 37.300000 ;
        RECT 372.120000 53.140000 373.320000 53.620000 ;
        RECT 372.120000 47.700000 373.320000 48.180000 ;
        RECT 372.120000 42.260000 373.320000 42.740000 ;
        RECT 372.120000 64.020000 373.320000 64.500000 ;
        RECT 372.120000 58.580000 373.320000 59.060000 ;
        RECT 372.120000 69.460000 373.320000 69.940000 ;
        RECT 417.120000 53.140000 418.320000 53.620000 ;
        RECT 417.120000 47.700000 418.320000 48.180000 ;
        RECT 417.120000 42.260000 418.320000 42.740000 ;
        RECT 417.120000 64.020000 418.320000 64.500000 ;
        RECT 417.120000 58.580000 418.320000 59.060000 ;
        RECT 417.120000 69.460000 418.320000 69.940000 ;
        RECT 282.120000 91.220000 283.320000 91.700000 ;
        RECT 282.120000 85.780000 283.320000 86.260000 ;
        RECT 282.120000 80.340000 283.320000 80.820000 ;
        RECT 282.120000 107.540000 283.320000 108.020000 ;
        RECT 282.120000 96.660000 283.320000 97.140000 ;
        RECT 282.120000 102.100000 283.320000 102.580000 ;
        RECT 327.120000 91.220000 328.320000 91.700000 ;
        RECT 327.120000 85.780000 328.320000 86.260000 ;
        RECT 327.120000 80.340000 328.320000 80.820000 ;
        RECT 327.120000 96.660000 328.320000 97.140000 ;
        RECT 327.120000 102.100000 328.320000 102.580000 ;
        RECT 327.120000 107.540000 328.320000 108.020000 ;
        RECT 282.120000 129.300000 283.320000 129.780000 ;
        RECT 282.120000 123.860000 283.320000 124.340000 ;
        RECT 282.120000 118.420000 283.320000 118.900000 ;
        RECT 282.120000 112.980000 283.320000 113.460000 ;
        RECT 282.120000 134.740000 283.320000 135.220000 ;
        RECT 282.120000 140.180000 283.320000 140.660000 ;
        RECT 282.120000 145.620000 283.320000 146.100000 ;
        RECT 327.120000 129.300000 328.320000 129.780000 ;
        RECT 327.120000 123.860000 328.320000 124.340000 ;
        RECT 327.120000 118.420000 328.320000 118.900000 ;
        RECT 327.120000 112.980000 328.320000 113.460000 ;
        RECT 327.120000 134.740000 328.320000 135.220000 ;
        RECT 327.120000 140.180000 328.320000 140.660000 ;
        RECT 327.120000 145.620000 328.320000 146.100000 ;
        RECT 372.120000 85.780000 373.320000 86.260000 ;
        RECT 372.120000 80.340000 373.320000 80.820000 ;
        RECT 372.120000 91.220000 373.320000 91.700000 ;
        RECT 372.120000 107.540000 373.320000 108.020000 ;
        RECT 372.120000 96.660000 373.320000 97.140000 ;
        RECT 372.120000 102.100000 373.320000 102.580000 ;
        RECT 417.120000 85.780000 418.320000 86.260000 ;
        RECT 417.120000 80.340000 418.320000 80.820000 ;
        RECT 417.120000 91.220000 418.320000 91.700000 ;
        RECT 417.120000 96.660000 418.320000 97.140000 ;
        RECT 417.120000 102.100000 418.320000 102.580000 ;
        RECT 417.120000 107.540000 418.320000 108.020000 ;
        RECT 372.120000 129.300000 373.320000 129.780000 ;
        RECT 372.120000 123.860000 373.320000 124.340000 ;
        RECT 372.120000 118.420000 373.320000 118.900000 ;
        RECT 372.120000 112.980000 373.320000 113.460000 ;
        RECT 372.120000 134.740000 373.320000 135.220000 ;
        RECT 372.120000 140.180000 373.320000 140.660000 ;
        RECT 372.120000 145.620000 373.320000 146.100000 ;
        RECT 417.120000 129.300000 418.320000 129.780000 ;
        RECT 417.120000 123.860000 418.320000 124.340000 ;
        RECT 417.120000 118.420000 418.320000 118.900000 ;
        RECT 417.120000 112.980000 418.320000 113.460000 ;
        RECT 417.120000 134.740000 418.320000 135.220000 ;
        RECT 417.120000 140.180000 418.320000 140.660000 ;
        RECT 417.120000 145.620000 418.320000 146.100000 ;
        RECT 543.400000 74.900000 544.600000 75.380000 ;
        RECT 507.120000 74.900000 508.320000 75.380000 ;
        RECT 462.120000 74.900000 463.320000 75.380000 ;
        RECT 462.120000 31.380000 463.320000 31.860000 ;
        RECT 462.120000 9.620000 463.320000 10.100000 ;
        RECT 462.120000 15.060000 463.320000 15.540000 ;
        RECT 462.120000 20.500000 463.320000 20.980000 ;
        RECT 462.120000 25.940000 463.320000 26.420000 ;
        RECT 462.120000 36.820000 463.320000 37.300000 ;
        RECT 462.120000 69.460000 463.320000 69.940000 ;
        RECT 462.120000 64.020000 463.320000 64.500000 ;
        RECT 462.120000 42.260000 463.320000 42.740000 ;
        RECT 462.120000 47.700000 463.320000 48.180000 ;
        RECT 462.120000 53.140000 463.320000 53.620000 ;
        RECT 462.120000 58.580000 463.320000 59.060000 ;
        RECT 507.120000 9.620000 508.320000 10.100000 ;
        RECT 507.120000 15.060000 508.320000 15.540000 ;
        RECT 507.120000 20.500000 508.320000 20.980000 ;
        RECT 507.120000 25.940000 508.320000 26.420000 ;
        RECT 507.120000 31.380000 508.320000 31.860000 ;
        RECT 507.120000 36.820000 508.320000 37.300000 ;
        RECT 543.400000 15.060000 544.600000 15.540000 ;
        RECT 543.400000 9.620000 544.600000 10.100000 ;
        RECT 543.400000 36.820000 544.600000 37.300000 ;
        RECT 543.400000 31.380000 544.600000 31.860000 ;
        RECT 543.400000 25.940000 544.600000 26.420000 ;
        RECT 543.400000 20.500000 544.600000 20.980000 ;
        RECT 507.120000 42.260000 508.320000 42.740000 ;
        RECT 507.120000 47.700000 508.320000 48.180000 ;
        RECT 507.120000 53.140000 508.320000 53.620000 ;
        RECT 507.120000 69.460000 508.320000 69.940000 ;
        RECT 507.120000 64.020000 508.320000 64.500000 ;
        RECT 507.120000 58.580000 508.320000 59.060000 ;
        RECT 543.400000 53.140000 544.600000 53.620000 ;
        RECT 543.400000 47.700000 544.600000 48.180000 ;
        RECT 543.400000 42.260000 544.600000 42.740000 ;
        RECT 543.400000 69.460000 544.600000 69.940000 ;
        RECT 543.400000 64.020000 544.600000 64.500000 ;
        RECT 543.400000 58.580000 544.600000 59.060000 ;
        RECT 462.120000 102.100000 463.320000 102.580000 ;
        RECT 462.120000 96.660000 463.320000 97.140000 ;
        RECT 462.120000 91.220000 463.320000 91.700000 ;
        RECT 462.120000 85.780000 463.320000 86.260000 ;
        RECT 462.120000 80.340000 463.320000 80.820000 ;
        RECT 462.120000 107.540000 463.320000 108.020000 ;
        RECT 462.120000 145.620000 463.320000 146.100000 ;
        RECT 462.120000 140.180000 463.320000 140.660000 ;
        RECT 462.120000 134.740000 463.320000 135.220000 ;
        RECT 462.120000 112.980000 463.320000 113.460000 ;
        RECT 462.120000 118.420000 463.320000 118.900000 ;
        RECT 462.120000 123.860000 463.320000 124.340000 ;
        RECT 462.120000 129.300000 463.320000 129.780000 ;
        RECT 507.120000 91.220000 508.320000 91.700000 ;
        RECT 507.120000 85.780000 508.320000 86.260000 ;
        RECT 507.120000 80.340000 508.320000 80.820000 ;
        RECT 507.120000 102.100000 508.320000 102.580000 ;
        RECT 507.120000 96.660000 508.320000 97.140000 ;
        RECT 507.120000 107.540000 508.320000 108.020000 ;
        RECT 543.400000 91.220000 544.600000 91.700000 ;
        RECT 543.400000 85.780000 544.600000 86.260000 ;
        RECT 543.400000 80.340000 544.600000 80.820000 ;
        RECT 543.400000 107.540000 544.600000 108.020000 ;
        RECT 543.400000 102.100000 544.600000 102.580000 ;
        RECT 543.400000 96.660000 544.600000 97.140000 ;
        RECT 507.120000 112.980000 508.320000 113.460000 ;
        RECT 507.120000 118.420000 508.320000 118.900000 ;
        RECT 507.120000 123.860000 508.320000 124.340000 ;
        RECT 507.120000 129.300000 508.320000 129.780000 ;
        RECT 507.120000 145.620000 508.320000 146.100000 ;
        RECT 507.120000 140.180000 508.320000 140.660000 ;
        RECT 507.120000 134.740000 508.320000 135.220000 ;
        RECT 543.400000 129.300000 544.600000 129.780000 ;
        RECT 543.400000 123.860000 544.600000 124.340000 ;
        RECT 543.400000 118.420000 544.600000 118.900000 ;
        RECT 543.400000 112.980000 544.600000 113.460000 ;
        RECT 543.400000 145.620000 544.600000 146.100000 ;
        RECT 543.400000 140.180000 544.600000 140.660000 ;
        RECT 543.400000 134.740000 544.600000 135.220000 ;
        RECT 282.120000 156.500000 283.320000 156.980000 ;
        RECT 282.120000 151.060000 283.320000 151.540000 ;
        RECT 282.120000 161.940000 283.320000 162.420000 ;
        RECT 282.120000 167.380000 283.320000 167.860000 ;
        RECT 282.120000 178.260000 283.320000 178.740000 ;
        RECT 282.120000 172.820000 283.320000 173.300000 ;
        RECT 282.120000 183.700000 283.320000 184.180000 ;
        RECT 327.120000 156.500000 328.320000 156.980000 ;
        RECT 327.120000 151.060000 328.320000 151.540000 ;
        RECT 327.120000 161.940000 328.320000 162.420000 ;
        RECT 327.120000 167.380000 328.320000 167.860000 ;
        RECT 327.120000 172.820000 328.320000 173.300000 ;
        RECT 327.120000 178.260000 328.320000 178.740000 ;
        RECT 327.120000 183.700000 328.320000 184.180000 ;
        RECT 282.120000 205.460000 283.320000 205.940000 ;
        RECT 282.120000 200.020000 283.320000 200.500000 ;
        RECT 282.120000 194.580000 283.320000 195.060000 ;
        RECT 282.120000 189.140000 283.320000 189.620000 ;
        RECT 282.120000 210.900000 283.320000 211.380000 ;
        RECT 282.120000 216.340000 283.320000 216.820000 ;
        RECT 282.120000 221.780000 283.320000 222.260000 ;
        RECT 327.120000 205.460000 328.320000 205.940000 ;
        RECT 327.120000 200.020000 328.320000 200.500000 ;
        RECT 327.120000 194.580000 328.320000 195.060000 ;
        RECT 327.120000 189.140000 328.320000 189.620000 ;
        RECT 327.120000 210.900000 328.320000 211.380000 ;
        RECT 327.120000 216.340000 328.320000 216.820000 ;
        RECT 327.120000 221.780000 328.320000 222.260000 ;
        RECT 372.120000 161.940000 373.320000 162.420000 ;
        RECT 372.120000 156.500000 373.320000 156.980000 ;
        RECT 372.120000 151.060000 373.320000 151.540000 ;
        RECT 372.120000 167.380000 373.320000 167.860000 ;
        RECT 372.120000 178.260000 373.320000 178.740000 ;
        RECT 372.120000 172.820000 373.320000 173.300000 ;
        RECT 372.120000 183.700000 373.320000 184.180000 ;
        RECT 417.120000 156.500000 418.320000 156.980000 ;
        RECT 417.120000 151.060000 418.320000 151.540000 ;
        RECT 417.120000 161.940000 418.320000 162.420000 ;
        RECT 417.120000 167.380000 418.320000 167.860000 ;
        RECT 417.120000 172.820000 418.320000 173.300000 ;
        RECT 417.120000 178.260000 418.320000 178.740000 ;
        RECT 417.120000 183.700000 418.320000 184.180000 ;
        RECT 372.120000 205.460000 373.320000 205.940000 ;
        RECT 372.120000 200.020000 373.320000 200.500000 ;
        RECT 372.120000 194.580000 373.320000 195.060000 ;
        RECT 372.120000 189.140000 373.320000 189.620000 ;
        RECT 372.120000 210.900000 373.320000 211.380000 ;
        RECT 372.120000 216.340000 373.320000 216.820000 ;
        RECT 372.120000 221.780000 373.320000 222.260000 ;
        RECT 417.120000 205.460000 418.320000 205.940000 ;
        RECT 417.120000 200.020000 418.320000 200.500000 ;
        RECT 417.120000 194.580000 418.320000 195.060000 ;
        RECT 417.120000 189.140000 418.320000 189.620000 ;
        RECT 417.120000 210.900000 418.320000 211.380000 ;
        RECT 417.120000 216.340000 418.320000 216.820000 ;
        RECT 417.120000 221.780000 418.320000 222.260000 ;
        RECT 282.120000 243.540000 283.320000 244.020000 ;
        RECT 282.120000 238.100000 283.320000 238.580000 ;
        RECT 282.120000 232.660000 283.320000 233.140000 ;
        RECT 282.120000 227.220000 283.320000 227.700000 ;
        RECT 282.120000 254.420000 283.320000 254.900000 ;
        RECT 282.120000 248.980000 283.320000 249.460000 ;
        RECT 282.120000 259.860000 283.320000 260.340000 ;
        RECT 327.120000 243.540000 328.320000 244.020000 ;
        RECT 327.120000 238.100000 328.320000 238.580000 ;
        RECT 327.120000 232.660000 328.320000 233.140000 ;
        RECT 327.120000 227.220000 328.320000 227.700000 ;
        RECT 327.120000 248.980000 328.320000 249.460000 ;
        RECT 327.120000 254.420000 328.320000 254.900000 ;
        RECT 327.120000 259.860000 328.320000 260.340000 ;
        RECT 282.120000 276.180000 283.320000 276.660000 ;
        RECT 282.120000 270.740000 283.320000 271.220000 ;
        RECT 282.120000 265.300000 283.320000 265.780000 ;
        RECT 282.120000 287.060000 283.320000 287.540000 ;
        RECT 282.120000 281.620000 283.320000 282.100000 ;
        RECT 282.120000 292.500000 283.320000 292.980000 ;
        RECT 282.120000 297.940000 283.320000 298.420000 ;
        RECT 327.120000 276.180000 328.320000 276.660000 ;
        RECT 327.120000 270.740000 328.320000 271.220000 ;
        RECT 327.120000 265.300000 328.320000 265.780000 ;
        RECT 327.120000 287.060000 328.320000 287.540000 ;
        RECT 327.120000 281.620000 328.320000 282.100000 ;
        RECT 327.120000 292.500000 328.320000 292.980000 ;
        RECT 327.120000 297.940000 328.320000 298.420000 ;
        RECT 372.120000 243.540000 373.320000 244.020000 ;
        RECT 372.120000 232.660000 373.320000 233.140000 ;
        RECT 372.120000 227.220000 373.320000 227.700000 ;
        RECT 372.120000 238.100000 373.320000 238.580000 ;
        RECT 372.120000 254.420000 373.320000 254.900000 ;
        RECT 372.120000 248.980000 373.320000 249.460000 ;
        RECT 372.120000 259.860000 373.320000 260.340000 ;
        RECT 417.120000 243.540000 418.320000 244.020000 ;
        RECT 417.120000 232.660000 418.320000 233.140000 ;
        RECT 417.120000 227.220000 418.320000 227.700000 ;
        RECT 417.120000 238.100000 418.320000 238.580000 ;
        RECT 417.120000 248.980000 418.320000 249.460000 ;
        RECT 417.120000 254.420000 418.320000 254.900000 ;
        RECT 417.120000 259.860000 418.320000 260.340000 ;
        RECT 372.120000 276.180000 373.320000 276.660000 ;
        RECT 372.120000 270.740000 373.320000 271.220000 ;
        RECT 372.120000 265.300000 373.320000 265.780000 ;
        RECT 372.120000 287.060000 373.320000 287.540000 ;
        RECT 372.120000 281.620000 373.320000 282.100000 ;
        RECT 372.120000 292.500000 373.320000 292.980000 ;
        RECT 372.120000 297.940000 373.320000 298.420000 ;
        RECT 417.120000 276.180000 418.320000 276.660000 ;
        RECT 417.120000 270.740000 418.320000 271.220000 ;
        RECT 417.120000 265.300000 418.320000 265.780000 ;
        RECT 417.120000 287.060000 418.320000 287.540000 ;
        RECT 417.120000 281.620000 418.320000 282.100000 ;
        RECT 417.120000 292.500000 418.320000 292.980000 ;
        RECT 417.120000 297.940000 418.320000 298.420000 ;
        RECT 462.120000 178.260000 463.320000 178.740000 ;
        RECT 462.120000 151.060000 463.320000 151.540000 ;
        RECT 462.120000 156.500000 463.320000 156.980000 ;
        RECT 462.120000 161.940000 463.320000 162.420000 ;
        RECT 462.120000 167.380000 463.320000 167.860000 ;
        RECT 462.120000 172.820000 463.320000 173.300000 ;
        RECT 462.120000 183.700000 463.320000 184.180000 ;
        RECT 462.120000 221.780000 463.320000 222.260000 ;
        RECT 462.120000 216.340000 463.320000 216.820000 ;
        RECT 462.120000 210.900000 463.320000 211.380000 ;
        RECT 462.120000 205.460000 463.320000 205.940000 ;
        RECT 462.120000 189.140000 463.320000 189.620000 ;
        RECT 462.120000 194.580000 463.320000 195.060000 ;
        RECT 462.120000 200.020000 463.320000 200.500000 ;
        RECT 507.120000 151.060000 508.320000 151.540000 ;
        RECT 507.120000 156.500000 508.320000 156.980000 ;
        RECT 507.120000 161.940000 508.320000 162.420000 ;
        RECT 507.120000 167.380000 508.320000 167.860000 ;
        RECT 507.120000 172.820000 508.320000 173.300000 ;
        RECT 507.120000 178.260000 508.320000 178.740000 ;
        RECT 507.120000 183.700000 508.320000 184.180000 ;
        RECT 543.400000 167.380000 544.600000 167.860000 ;
        RECT 543.400000 161.940000 544.600000 162.420000 ;
        RECT 543.400000 156.500000 544.600000 156.980000 ;
        RECT 543.400000 151.060000 544.600000 151.540000 ;
        RECT 543.400000 183.700000 544.600000 184.180000 ;
        RECT 543.400000 178.260000 544.600000 178.740000 ;
        RECT 543.400000 172.820000 544.600000 173.300000 ;
        RECT 507.120000 205.460000 508.320000 205.940000 ;
        RECT 507.120000 189.140000 508.320000 189.620000 ;
        RECT 507.120000 194.580000 508.320000 195.060000 ;
        RECT 507.120000 200.020000 508.320000 200.500000 ;
        RECT 507.120000 221.780000 508.320000 222.260000 ;
        RECT 507.120000 216.340000 508.320000 216.820000 ;
        RECT 507.120000 210.900000 508.320000 211.380000 ;
        RECT 543.400000 205.460000 544.600000 205.940000 ;
        RECT 543.400000 200.020000 544.600000 200.500000 ;
        RECT 543.400000 194.580000 544.600000 195.060000 ;
        RECT 543.400000 189.140000 544.600000 189.620000 ;
        RECT 543.400000 221.780000 544.600000 222.260000 ;
        RECT 543.400000 216.340000 544.600000 216.820000 ;
        RECT 543.400000 210.900000 544.600000 211.380000 ;
        RECT 462.120000 248.980000 463.320000 249.460000 ;
        RECT 462.120000 243.540000 463.320000 244.020000 ;
        RECT 462.120000 238.100000 463.320000 238.580000 ;
        RECT 462.120000 232.660000 463.320000 233.140000 ;
        RECT 462.120000 227.220000 463.320000 227.700000 ;
        RECT 462.120000 254.420000 463.320000 254.900000 ;
        RECT 462.120000 259.860000 463.320000 260.340000 ;
        RECT 462.120000 297.940000 463.320000 298.420000 ;
        RECT 462.120000 292.500000 463.320000 292.980000 ;
        RECT 462.120000 287.060000 463.320000 287.540000 ;
        RECT 462.120000 281.620000 463.320000 282.100000 ;
        RECT 462.120000 265.300000 463.320000 265.780000 ;
        RECT 462.120000 270.740000 463.320000 271.220000 ;
        RECT 462.120000 276.180000 463.320000 276.660000 ;
        RECT 507.120000 243.540000 508.320000 244.020000 ;
        RECT 507.120000 238.100000 508.320000 238.580000 ;
        RECT 507.120000 232.660000 508.320000 233.140000 ;
        RECT 507.120000 227.220000 508.320000 227.700000 ;
        RECT 507.120000 248.980000 508.320000 249.460000 ;
        RECT 507.120000 254.420000 508.320000 254.900000 ;
        RECT 507.120000 259.860000 508.320000 260.340000 ;
        RECT 543.400000 243.540000 544.600000 244.020000 ;
        RECT 543.400000 238.100000 544.600000 238.580000 ;
        RECT 543.400000 232.660000 544.600000 233.140000 ;
        RECT 543.400000 227.220000 544.600000 227.700000 ;
        RECT 543.400000 259.860000 544.600000 260.340000 ;
        RECT 543.400000 254.420000 544.600000 254.900000 ;
        RECT 543.400000 248.980000 544.600000 249.460000 ;
        RECT 507.120000 265.300000 508.320000 265.780000 ;
        RECT 507.120000 270.740000 508.320000 271.220000 ;
        RECT 507.120000 276.180000 508.320000 276.660000 ;
        RECT 507.120000 297.940000 508.320000 298.420000 ;
        RECT 507.120000 292.500000 508.320000 292.980000 ;
        RECT 507.120000 287.060000 508.320000 287.540000 ;
        RECT 507.120000 281.620000 508.320000 282.100000 ;
        RECT 543.400000 276.180000 544.600000 276.660000 ;
        RECT 543.400000 270.740000 544.600000 271.220000 ;
        RECT 543.400000 265.300000 544.600000 265.780000 ;
        RECT 543.400000 297.940000 544.600000 298.420000 ;
        RECT 543.400000 292.500000 544.600000 292.980000 ;
        RECT 543.400000 287.060000 544.600000 287.540000 ;
        RECT 543.400000 281.620000 544.600000 282.100000 ;
        RECT 12.120000 308.820000 13.320000 309.300000 ;
        RECT 12.120000 303.380000 13.320000 303.860000 ;
        RECT 12.120000 314.260000 13.320000 314.740000 ;
        RECT 12.120000 319.700000 13.320000 320.180000 ;
        RECT 12.120000 325.140000 13.320000 325.620000 ;
        RECT 12.120000 330.580000 13.320000 331.060000 ;
        RECT 12.120000 336.020000 13.320000 336.500000 ;
        RECT 5.560000 308.820000 6.760000 309.300000 ;
        RECT 5.560000 303.380000 6.760000 303.860000 ;
        RECT 5.560000 314.260000 6.760000 314.740000 ;
        RECT 5.560000 319.700000 6.760000 320.180000 ;
        RECT 5.560000 325.140000 6.760000 325.620000 ;
        RECT 5.560000 336.020000 6.760000 336.500000 ;
        RECT 5.560000 330.580000 6.760000 331.060000 ;
        RECT 12.120000 374.100000 13.320000 374.580000 ;
        RECT 12.120000 368.660000 13.320000 369.140000 ;
        RECT 12.120000 363.220000 13.320000 363.700000 ;
        RECT 12.120000 357.780000 13.320000 358.260000 ;
        RECT 12.120000 341.460000 13.320000 341.940000 ;
        RECT 12.120000 346.900000 13.320000 347.380000 ;
        RECT 12.120000 352.340000 13.320000 352.820000 ;
        RECT 5.560000 341.460000 6.760000 341.940000 ;
        RECT 5.560000 346.900000 6.760000 347.380000 ;
        RECT 5.560000 352.340000 6.760000 352.820000 ;
        RECT 5.560000 357.780000 6.760000 358.260000 ;
        RECT 5.560000 363.220000 6.760000 363.700000 ;
        RECT 5.560000 374.100000 6.760000 374.580000 ;
        RECT 5.560000 368.660000 6.760000 369.140000 ;
        RECT 57.120000 308.820000 58.320000 309.300000 ;
        RECT 57.120000 303.380000 58.320000 303.860000 ;
        RECT 57.120000 314.260000 58.320000 314.740000 ;
        RECT 57.120000 330.580000 58.320000 331.060000 ;
        RECT 57.120000 319.700000 58.320000 320.180000 ;
        RECT 57.120000 325.140000 58.320000 325.620000 ;
        RECT 57.120000 336.020000 58.320000 336.500000 ;
        RECT 102.120000 308.820000 103.320000 309.300000 ;
        RECT 102.120000 303.380000 103.320000 303.860000 ;
        RECT 102.120000 314.260000 103.320000 314.740000 ;
        RECT 102.120000 319.700000 103.320000 320.180000 ;
        RECT 102.120000 325.140000 103.320000 325.620000 ;
        RECT 102.120000 330.580000 103.320000 331.060000 ;
        RECT 102.120000 336.020000 103.320000 336.500000 ;
        RECT 57.120000 352.340000 58.320000 352.820000 ;
        RECT 57.120000 346.900000 58.320000 347.380000 ;
        RECT 57.120000 341.460000 58.320000 341.940000 ;
        RECT 57.120000 363.220000 58.320000 363.700000 ;
        RECT 57.120000 357.780000 58.320000 358.260000 ;
        RECT 57.120000 368.660000 58.320000 369.140000 ;
        RECT 57.120000 374.100000 58.320000 374.580000 ;
        RECT 102.120000 352.340000 103.320000 352.820000 ;
        RECT 102.120000 346.900000 103.320000 347.380000 ;
        RECT 102.120000 341.460000 103.320000 341.940000 ;
        RECT 102.120000 363.220000 103.320000 363.700000 ;
        RECT 102.120000 357.780000 103.320000 358.260000 ;
        RECT 102.120000 368.660000 103.320000 369.140000 ;
        RECT 102.120000 374.100000 103.320000 374.580000 ;
        RECT 5.560000 412.180000 6.760000 412.660000 ;
        RECT 12.120000 412.180000 13.320000 412.660000 ;
        RECT 12.120000 395.860000 13.320000 396.340000 ;
        RECT 12.120000 390.420000 13.320000 390.900000 ;
        RECT 12.120000 384.980000 13.320000 385.460000 ;
        RECT 12.120000 379.540000 13.320000 380.020000 ;
        RECT 12.120000 401.300000 13.320000 401.780000 ;
        RECT 12.120000 406.740000 13.320000 407.220000 ;
        RECT 5.560000 379.540000 6.760000 380.020000 ;
        RECT 5.560000 384.980000 6.760000 385.460000 ;
        RECT 5.560000 390.420000 6.760000 390.900000 ;
        RECT 5.560000 395.860000 6.760000 396.340000 ;
        RECT 5.560000 401.300000 6.760000 401.780000 ;
        RECT 5.560000 406.740000 6.760000 407.220000 ;
        RECT 12.120000 444.820000 13.320000 445.300000 ;
        RECT 12.120000 439.380000 13.320000 439.860000 ;
        RECT 12.120000 433.940000 13.320000 434.420000 ;
        RECT 12.120000 417.620000 13.320000 418.100000 ;
        RECT 12.120000 423.060000 13.320000 423.540000 ;
        RECT 12.120000 428.500000 13.320000 428.980000 ;
        RECT 5.560000 417.620000 6.760000 418.100000 ;
        RECT 5.560000 423.060000 6.760000 423.540000 ;
        RECT 5.560000 428.500000 6.760000 428.980000 ;
        RECT 5.560000 433.940000 6.760000 434.420000 ;
        RECT 5.560000 439.380000 6.760000 439.860000 ;
        RECT 5.560000 444.820000 6.760000 445.300000 ;
        RECT 102.120000 412.180000 103.320000 412.660000 ;
        RECT 57.120000 412.180000 58.320000 412.660000 ;
        RECT 57.120000 390.420000 58.320000 390.900000 ;
        RECT 57.120000 384.980000 58.320000 385.460000 ;
        RECT 57.120000 379.540000 58.320000 380.020000 ;
        RECT 57.120000 406.740000 58.320000 407.220000 ;
        RECT 57.120000 395.860000 58.320000 396.340000 ;
        RECT 57.120000 401.300000 58.320000 401.780000 ;
        RECT 102.120000 390.420000 103.320000 390.900000 ;
        RECT 102.120000 384.980000 103.320000 385.460000 ;
        RECT 102.120000 379.540000 103.320000 380.020000 ;
        RECT 102.120000 395.860000 103.320000 396.340000 ;
        RECT 102.120000 401.300000 103.320000 401.780000 ;
        RECT 102.120000 406.740000 103.320000 407.220000 ;
        RECT 57.120000 428.500000 58.320000 428.980000 ;
        RECT 57.120000 423.060000 58.320000 423.540000 ;
        RECT 57.120000 417.620000 58.320000 418.100000 ;
        RECT 57.120000 439.380000 58.320000 439.860000 ;
        RECT 57.120000 433.940000 58.320000 434.420000 ;
        RECT 57.120000 444.820000 58.320000 445.300000 ;
        RECT 102.120000 428.500000 103.320000 428.980000 ;
        RECT 102.120000 423.060000 103.320000 423.540000 ;
        RECT 102.120000 417.620000 103.320000 418.100000 ;
        RECT 102.120000 439.380000 103.320000 439.860000 ;
        RECT 102.120000 433.940000 103.320000 434.420000 ;
        RECT 102.120000 444.820000 103.320000 445.300000 ;
        RECT 147.120000 303.380000 148.320000 303.860000 ;
        RECT 147.120000 308.820000 148.320000 309.300000 ;
        RECT 147.120000 314.260000 148.320000 314.740000 ;
        RECT 147.120000 330.580000 148.320000 331.060000 ;
        RECT 147.120000 319.700000 148.320000 320.180000 ;
        RECT 147.120000 325.140000 148.320000 325.620000 ;
        RECT 147.120000 336.020000 148.320000 336.500000 ;
        RECT 192.120000 303.380000 193.320000 303.860000 ;
        RECT 192.120000 308.820000 193.320000 309.300000 ;
        RECT 192.120000 314.260000 193.320000 314.740000 ;
        RECT 192.120000 319.700000 193.320000 320.180000 ;
        RECT 192.120000 325.140000 193.320000 325.620000 ;
        RECT 192.120000 330.580000 193.320000 331.060000 ;
        RECT 192.120000 336.020000 193.320000 336.500000 ;
        RECT 147.120000 352.340000 148.320000 352.820000 ;
        RECT 147.120000 346.900000 148.320000 347.380000 ;
        RECT 147.120000 341.460000 148.320000 341.940000 ;
        RECT 147.120000 363.220000 148.320000 363.700000 ;
        RECT 147.120000 357.780000 148.320000 358.260000 ;
        RECT 147.120000 368.660000 148.320000 369.140000 ;
        RECT 147.120000 374.100000 148.320000 374.580000 ;
        RECT 192.120000 352.340000 193.320000 352.820000 ;
        RECT 192.120000 346.900000 193.320000 347.380000 ;
        RECT 192.120000 341.460000 193.320000 341.940000 ;
        RECT 192.120000 363.220000 193.320000 363.700000 ;
        RECT 192.120000 357.780000 193.320000 358.260000 ;
        RECT 192.120000 368.660000 193.320000 369.140000 ;
        RECT 192.120000 374.100000 193.320000 374.580000 ;
        RECT 237.120000 308.820000 238.320000 309.300000 ;
        RECT 237.120000 303.380000 238.320000 303.860000 ;
        RECT 237.120000 314.260000 238.320000 314.740000 ;
        RECT 237.120000 319.700000 238.320000 320.180000 ;
        RECT 237.120000 325.140000 238.320000 325.620000 ;
        RECT 237.120000 330.580000 238.320000 331.060000 ;
        RECT 237.120000 336.020000 238.320000 336.500000 ;
        RECT 237.120000 374.100000 238.320000 374.580000 ;
        RECT 237.120000 368.660000 238.320000 369.140000 ;
        RECT 237.120000 363.220000 238.320000 363.700000 ;
        RECT 237.120000 357.780000 238.320000 358.260000 ;
        RECT 237.120000 341.460000 238.320000 341.940000 ;
        RECT 237.120000 346.900000 238.320000 347.380000 ;
        RECT 237.120000 352.340000 238.320000 352.820000 ;
        RECT 192.120000 412.180000 193.320000 412.660000 ;
        RECT 147.120000 412.180000 148.320000 412.660000 ;
        RECT 147.120000 390.420000 148.320000 390.900000 ;
        RECT 147.120000 384.980000 148.320000 385.460000 ;
        RECT 147.120000 379.540000 148.320000 380.020000 ;
        RECT 147.120000 406.740000 148.320000 407.220000 ;
        RECT 147.120000 395.860000 148.320000 396.340000 ;
        RECT 147.120000 401.300000 148.320000 401.780000 ;
        RECT 192.120000 390.420000 193.320000 390.900000 ;
        RECT 192.120000 384.980000 193.320000 385.460000 ;
        RECT 192.120000 379.540000 193.320000 380.020000 ;
        RECT 192.120000 395.860000 193.320000 396.340000 ;
        RECT 192.120000 401.300000 193.320000 401.780000 ;
        RECT 192.120000 406.740000 193.320000 407.220000 ;
        RECT 147.120000 428.500000 148.320000 428.980000 ;
        RECT 147.120000 423.060000 148.320000 423.540000 ;
        RECT 147.120000 417.620000 148.320000 418.100000 ;
        RECT 147.120000 439.380000 148.320000 439.860000 ;
        RECT 147.120000 433.940000 148.320000 434.420000 ;
        RECT 147.120000 444.820000 148.320000 445.300000 ;
        RECT 192.120000 428.500000 193.320000 428.980000 ;
        RECT 192.120000 423.060000 193.320000 423.540000 ;
        RECT 192.120000 417.620000 193.320000 418.100000 ;
        RECT 192.120000 439.380000 193.320000 439.860000 ;
        RECT 192.120000 433.940000 193.320000 434.420000 ;
        RECT 192.120000 444.820000 193.320000 445.300000 ;
        RECT 237.120000 412.180000 238.320000 412.660000 ;
        RECT 237.120000 395.860000 238.320000 396.340000 ;
        RECT 237.120000 390.420000 238.320000 390.900000 ;
        RECT 237.120000 384.980000 238.320000 385.460000 ;
        RECT 237.120000 379.540000 238.320000 380.020000 ;
        RECT 237.120000 401.300000 238.320000 401.780000 ;
        RECT 237.120000 406.740000 238.320000 407.220000 ;
        RECT 237.120000 444.820000 238.320000 445.300000 ;
        RECT 237.120000 439.380000 238.320000 439.860000 ;
        RECT 237.120000 433.940000 238.320000 434.420000 ;
        RECT 237.120000 417.620000 238.320000 418.100000 ;
        RECT 237.120000 423.060000 238.320000 423.540000 ;
        RECT 237.120000 428.500000 238.320000 428.980000 ;
        RECT 12.120000 466.580000 13.320000 467.060000 ;
        RECT 12.120000 450.260000 13.320000 450.740000 ;
        RECT 12.120000 455.700000 13.320000 456.180000 ;
        RECT 12.120000 461.140000 13.320000 461.620000 ;
        RECT 12.120000 472.020000 13.320000 472.500000 ;
        RECT 12.120000 477.460000 13.320000 477.940000 ;
        RECT 12.120000 482.900000 13.320000 483.380000 ;
        RECT 5.560000 450.260000 6.760000 450.740000 ;
        RECT 5.560000 455.700000 6.760000 456.180000 ;
        RECT 5.560000 461.140000 6.760000 461.620000 ;
        RECT 5.560000 466.580000 6.760000 467.060000 ;
        RECT 5.560000 477.460000 6.760000 477.940000 ;
        RECT 5.560000 472.020000 6.760000 472.500000 ;
        RECT 5.560000 482.900000 6.760000 483.380000 ;
        RECT 12.120000 520.980000 13.320000 521.460000 ;
        RECT 12.120000 515.540000 13.320000 516.020000 ;
        RECT 12.120000 510.100000 13.320000 510.580000 ;
        RECT 12.120000 504.660000 13.320000 505.140000 ;
        RECT 12.120000 488.340000 13.320000 488.820000 ;
        RECT 12.120000 493.780000 13.320000 494.260000 ;
        RECT 12.120000 499.220000 13.320000 499.700000 ;
        RECT 5.560000 488.340000 6.760000 488.820000 ;
        RECT 5.560000 493.780000 6.760000 494.260000 ;
        RECT 5.560000 499.220000 6.760000 499.700000 ;
        RECT 5.560000 504.660000 6.760000 505.140000 ;
        RECT 5.560000 510.100000 6.760000 510.580000 ;
        RECT 5.560000 520.980000 6.760000 521.460000 ;
        RECT 5.560000 515.540000 6.760000 516.020000 ;
        RECT 57.120000 450.260000 58.320000 450.740000 ;
        RECT 57.120000 455.700000 58.320000 456.180000 ;
        RECT 57.120000 461.140000 58.320000 461.620000 ;
        RECT 57.120000 466.580000 58.320000 467.060000 ;
        RECT 57.120000 477.460000 58.320000 477.940000 ;
        RECT 57.120000 472.020000 58.320000 472.500000 ;
        RECT 57.120000 482.900000 58.320000 483.380000 ;
        RECT 102.120000 461.140000 103.320000 461.620000 ;
        RECT 102.120000 450.260000 103.320000 450.740000 ;
        RECT 102.120000 455.700000 103.320000 456.180000 ;
        RECT 102.120000 466.580000 103.320000 467.060000 ;
        RECT 102.120000 472.020000 103.320000 472.500000 ;
        RECT 102.120000 477.460000 103.320000 477.940000 ;
        RECT 102.120000 482.900000 103.320000 483.380000 ;
        RECT 57.120000 504.660000 58.320000 505.140000 ;
        RECT 57.120000 499.220000 58.320000 499.700000 ;
        RECT 57.120000 493.780000 58.320000 494.260000 ;
        RECT 57.120000 488.340000 58.320000 488.820000 ;
        RECT 57.120000 510.100000 58.320000 510.580000 ;
        RECT 57.120000 515.540000 58.320000 516.020000 ;
        RECT 57.120000 520.980000 58.320000 521.460000 ;
        RECT 102.120000 504.660000 103.320000 505.140000 ;
        RECT 102.120000 499.220000 103.320000 499.700000 ;
        RECT 102.120000 493.780000 103.320000 494.260000 ;
        RECT 102.120000 488.340000 103.320000 488.820000 ;
        RECT 102.120000 510.100000 103.320000 510.580000 ;
        RECT 102.120000 515.540000 103.320000 516.020000 ;
        RECT 102.120000 520.980000 103.320000 521.460000 ;
        RECT 12.120000 537.300000 13.320000 537.780000 ;
        RECT 12.120000 531.860000 13.320000 532.340000 ;
        RECT 12.120000 526.420000 13.320000 526.900000 ;
        RECT 12.120000 542.740000 13.320000 543.220000 ;
        RECT 12.120000 548.180000 13.320000 548.660000 ;
        RECT 12.120000 553.620000 13.320000 554.100000 ;
        RECT 12.120000 559.060000 13.320000 559.540000 ;
        RECT 5.560000 526.420000 6.760000 526.900000 ;
        RECT 5.560000 531.860000 6.760000 532.340000 ;
        RECT 5.560000 537.300000 6.760000 537.780000 ;
        RECT 5.560000 542.740000 6.760000 543.220000 ;
        RECT 5.560000 548.180000 6.760000 548.660000 ;
        RECT 5.560000 559.060000 6.760000 559.540000 ;
        RECT 5.560000 553.620000 6.760000 554.100000 ;
        RECT 12.120000 586.260000 13.320000 586.740000 ;
        RECT 12.120000 580.820000 13.320000 581.300000 ;
        RECT 12.120000 575.380000 13.320000 575.860000 ;
        RECT 12.120000 564.500000 13.320000 564.980000 ;
        RECT 12.120000 569.940000 13.320000 570.420000 ;
        RECT 5.560000 580.820000 6.760000 581.300000 ;
        RECT 5.560000 564.500000 6.760000 564.980000 ;
        RECT 5.560000 569.940000 6.760000 570.420000 ;
        RECT 5.560000 575.380000 6.760000 575.860000 ;
        RECT 5.560000 586.260000 6.760000 586.740000 ;
        RECT 57.120000 537.300000 58.320000 537.780000 ;
        RECT 57.120000 531.860000 58.320000 532.340000 ;
        RECT 57.120000 526.420000 58.320000 526.900000 ;
        RECT 57.120000 542.740000 58.320000 543.220000 ;
        RECT 57.120000 548.180000 58.320000 548.660000 ;
        RECT 57.120000 553.620000 58.320000 554.100000 ;
        RECT 57.120000 559.060000 58.320000 559.540000 ;
        RECT 102.120000 531.860000 103.320000 532.340000 ;
        RECT 102.120000 526.420000 103.320000 526.900000 ;
        RECT 102.120000 537.300000 103.320000 537.780000 ;
        RECT 102.120000 542.740000 103.320000 543.220000 ;
        RECT 102.120000 548.180000 103.320000 548.660000 ;
        RECT 102.120000 553.620000 103.320000 554.100000 ;
        RECT 102.120000 559.060000 103.320000 559.540000 ;
        RECT 57.120000 580.820000 58.320000 581.300000 ;
        RECT 57.120000 575.380000 58.320000 575.860000 ;
        RECT 57.120000 569.940000 58.320000 570.420000 ;
        RECT 57.120000 564.500000 58.320000 564.980000 ;
        RECT 57.120000 586.260000 58.320000 586.740000 ;
        RECT 102.120000 580.820000 103.320000 581.300000 ;
        RECT 102.120000 575.380000 103.320000 575.860000 ;
        RECT 102.120000 569.940000 103.320000 570.420000 ;
        RECT 102.120000 564.500000 103.320000 564.980000 ;
        RECT 102.120000 586.260000 103.320000 586.740000 ;
        RECT 147.120000 450.260000 148.320000 450.740000 ;
        RECT 147.120000 455.700000 148.320000 456.180000 ;
        RECT 147.120000 461.140000 148.320000 461.620000 ;
        RECT 147.120000 466.580000 148.320000 467.060000 ;
        RECT 147.120000 477.460000 148.320000 477.940000 ;
        RECT 147.120000 472.020000 148.320000 472.500000 ;
        RECT 147.120000 482.900000 148.320000 483.380000 ;
        RECT 192.120000 461.140000 193.320000 461.620000 ;
        RECT 192.120000 450.260000 193.320000 450.740000 ;
        RECT 192.120000 455.700000 193.320000 456.180000 ;
        RECT 192.120000 466.580000 193.320000 467.060000 ;
        RECT 192.120000 472.020000 193.320000 472.500000 ;
        RECT 192.120000 477.460000 193.320000 477.940000 ;
        RECT 192.120000 482.900000 193.320000 483.380000 ;
        RECT 147.120000 504.660000 148.320000 505.140000 ;
        RECT 147.120000 499.220000 148.320000 499.700000 ;
        RECT 147.120000 493.780000 148.320000 494.260000 ;
        RECT 147.120000 488.340000 148.320000 488.820000 ;
        RECT 147.120000 510.100000 148.320000 510.580000 ;
        RECT 147.120000 515.540000 148.320000 516.020000 ;
        RECT 147.120000 520.980000 148.320000 521.460000 ;
        RECT 192.120000 504.660000 193.320000 505.140000 ;
        RECT 192.120000 499.220000 193.320000 499.700000 ;
        RECT 192.120000 493.780000 193.320000 494.260000 ;
        RECT 192.120000 488.340000 193.320000 488.820000 ;
        RECT 192.120000 510.100000 193.320000 510.580000 ;
        RECT 192.120000 515.540000 193.320000 516.020000 ;
        RECT 192.120000 520.980000 193.320000 521.460000 ;
        RECT 237.120000 466.580000 238.320000 467.060000 ;
        RECT 237.120000 450.260000 238.320000 450.740000 ;
        RECT 237.120000 455.700000 238.320000 456.180000 ;
        RECT 237.120000 461.140000 238.320000 461.620000 ;
        RECT 237.120000 472.020000 238.320000 472.500000 ;
        RECT 237.120000 477.460000 238.320000 477.940000 ;
        RECT 237.120000 482.900000 238.320000 483.380000 ;
        RECT 237.120000 520.980000 238.320000 521.460000 ;
        RECT 237.120000 515.540000 238.320000 516.020000 ;
        RECT 237.120000 510.100000 238.320000 510.580000 ;
        RECT 237.120000 504.660000 238.320000 505.140000 ;
        RECT 237.120000 488.340000 238.320000 488.820000 ;
        RECT 237.120000 493.780000 238.320000 494.260000 ;
        RECT 237.120000 499.220000 238.320000 499.700000 ;
        RECT 147.120000 537.300000 148.320000 537.780000 ;
        RECT 147.120000 531.860000 148.320000 532.340000 ;
        RECT 147.120000 526.420000 148.320000 526.900000 ;
        RECT 147.120000 542.740000 148.320000 543.220000 ;
        RECT 147.120000 548.180000 148.320000 548.660000 ;
        RECT 147.120000 553.620000 148.320000 554.100000 ;
        RECT 147.120000 559.060000 148.320000 559.540000 ;
        RECT 192.120000 531.860000 193.320000 532.340000 ;
        RECT 192.120000 526.420000 193.320000 526.900000 ;
        RECT 192.120000 537.300000 193.320000 537.780000 ;
        RECT 192.120000 542.740000 193.320000 543.220000 ;
        RECT 192.120000 548.180000 193.320000 548.660000 ;
        RECT 192.120000 553.620000 193.320000 554.100000 ;
        RECT 192.120000 559.060000 193.320000 559.540000 ;
        RECT 147.120000 580.820000 148.320000 581.300000 ;
        RECT 147.120000 575.380000 148.320000 575.860000 ;
        RECT 147.120000 569.940000 148.320000 570.420000 ;
        RECT 147.120000 564.500000 148.320000 564.980000 ;
        RECT 147.120000 586.260000 148.320000 586.740000 ;
        RECT 192.120000 580.820000 193.320000 581.300000 ;
        RECT 192.120000 575.380000 193.320000 575.860000 ;
        RECT 192.120000 569.940000 193.320000 570.420000 ;
        RECT 192.120000 564.500000 193.320000 564.980000 ;
        RECT 192.120000 586.260000 193.320000 586.740000 ;
        RECT 237.120000 537.300000 238.320000 537.780000 ;
        RECT 237.120000 531.860000 238.320000 532.340000 ;
        RECT 237.120000 526.420000 238.320000 526.900000 ;
        RECT 237.120000 542.740000 238.320000 543.220000 ;
        RECT 237.120000 548.180000 238.320000 548.660000 ;
        RECT 237.120000 553.620000 238.320000 554.100000 ;
        RECT 237.120000 559.060000 238.320000 559.540000 ;
        RECT 237.120000 586.260000 238.320000 586.740000 ;
        RECT 237.120000 580.820000 238.320000 581.300000 ;
        RECT 237.120000 564.500000 238.320000 564.980000 ;
        RECT 237.120000 569.940000 238.320000 570.420000 ;
        RECT 237.120000 575.380000 238.320000 575.860000 ;
        RECT 282.120000 308.820000 283.320000 309.300000 ;
        RECT 282.120000 303.380000 283.320000 303.860000 ;
        RECT 282.120000 314.260000 283.320000 314.740000 ;
        RECT 282.120000 330.580000 283.320000 331.060000 ;
        RECT 282.120000 319.700000 283.320000 320.180000 ;
        RECT 282.120000 325.140000 283.320000 325.620000 ;
        RECT 282.120000 336.020000 283.320000 336.500000 ;
        RECT 327.120000 308.820000 328.320000 309.300000 ;
        RECT 327.120000 303.380000 328.320000 303.860000 ;
        RECT 327.120000 314.260000 328.320000 314.740000 ;
        RECT 327.120000 319.700000 328.320000 320.180000 ;
        RECT 327.120000 325.140000 328.320000 325.620000 ;
        RECT 327.120000 330.580000 328.320000 331.060000 ;
        RECT 327.120000 336.020000 328.320000 336.500000 ;
        RECT 282.120000 352.340000 283.320000 352.820000 ;
        RECT 282.120000 346.900000 283.320000 347.380000 ;
        RECT 282.120000 341.460000 283.320000 341.940000 ;
        RECT 282.120000 363.220000 283.320000 363.700000 ;
        RECT 282.120000 357.780000 283.320000 358.260000 ;
        RECT 282.120000 368.660000 283.320000 369.140000 ;
        RECT 282.120000 374.100000 283.320000 374.580000 ;
        RECT 327.120000 352.340000 328.320000 352.820000 ;
        RECT 327.120000 346.900000 328.320000 347.380000 ;
        RECT 327.120000 341.460000 328.320000 341.940000 ;
        RECT 327.120000 363.220000 328.320000 363.700000 ;
        RECT 327.120000 357.780000 328.320000 358.260000 ;
        RECT 327.120000 368.660000 328.320000 369.140000 ;
        RECT 327.120000 374.100000 328.320000 374.580000 ;
        RECT 372.120000 314.260000 373.320000 314.740000 ;
        RECT 372.120000 308.820000 373.320000 309.300000 ;
        RECT 372.120000 303.380000 373.320000 303.860000 ;
        RECT 372.120000 330.580000 373.320000 331.060000 ;
        RECT 372.120000 319.700000 373.320000 320.180000 ;
        RECT 372.120000 325.140000 373.320000 325.620000 ;
        RECT 372.120000 336.020000 373.320000 336.500000 ;
        RECT 417.120000 308.820000 418.320000 309.300000 ;
        RECT 417.120000 303.380000 418.320000 303.860000 ;
        RECT 417.120000 314.260000 418.320000 314.740000 ;
        RECT 417.120000 319.700000 418.320000 320.180000 ;
        RECT 417.120000 325.140000 418.320000 325.620000 ;
        RECT 417.120000 330.580000 418.320000 331.060000 ;
        RECT 417.120000 336.020000 418.320000 336.500000 ;
        RECT 372.120000 352.340000 373.320000 352.820000 ;
        RECT 372.120000 346.900000 373.320000 347.380000 ;
        RECT 372.120000 341.460000 373.320000 341.940000 ;
        RECT 372.120000 363.220000 373.320000 363.700000 ;
        RECT 372.120000 357.780000 373.320000 358.260000 ;
        RECT 372.120000 368.660000 373.320000 369.140000 ;
        RECT 372.120000 374.100000 373.320000 374.580000 ;
        RECT 417.120000 352.340000 418.320000 352.820000 ;
        RECT 417.120000 346.900000 418.320000 347.380000 ;
        RECT 417.120000 341.460000 418.320000 341.940000 ;
        RECT 417.120000 363.220000 418.320000 363.700000 ;
        RECT 417.120000 357.780000 418.320000 358.260000 ;
        RECT 417.120000 368.660000 418.320000 369.140000 ;
        RECT 417.120000 374.100000 418.320000 374.580000 ;
        RECT 327.120000 412.180000 328.320000 412.660000 ;
        RECT 282.120000 412.180000 283.320000 412.660000 ;
        RECT 282.120000 390.420000 283.320000 390.900000 ;
        RECT 282.120000 384.980000 283.320000 385.460000 ;
        RECT 282.120000 379.540000 283.320000 380.020000 ;
        RECT 282.120000 406.740000 283.320000 407.220000 ;
        RECT 282.120000 395.860000 283.320000 396.340000 ;
        RECT 282.120000 401.300000 283.320000 401.780000 ;
        RECT 327.120000 390.420000 328.320000 390.900000 ;
        RECT 327.120000 384.980000 328.320000 385.460000 ;
        RECT 327.120000 379.540000 328.320000 380.020000 ;
        RECT 327.120000 395.860000 328.320000 396.340000 ;
        RECT 327.120000 401.300000 328.320000 401.780000 ;
        RECT 327.120000 406.740000 328.320000 407.220000 ;
        RECT 282.120000 428.500000 283.320000 428.980000 ;
        RECT 282.120000 423.060000 283.320000 423.540000 ;
        RECT 282.120000 417.620000 283.320000 418.100000 ;
        RECT 282.120000 439.380000 283.320000 439.860000 ;
        RECT 282.120000 433.940000 283.320000 434.420000 ;
        RECT 282.120000 444.820000 283.320000 445.300000 ;
        RECT 327.120000 428.500000 328.320000 428.980000 ;
        RECT 327.120000 423.060000 328.320000 423.540000 ;
        RECT 327.120000 417.620000 328.320000 418.100000 ;
        RECT 327.120000 439.380000 328.320000 439.860000 ;
        RECT 327.120000 433.940000 328.320000 434.420000 ;
        RECT 327.120000 444.820000 328.320000 445.300000 ;
        RECT 417.120000 412.180000 418.320000 412.660000 ;
        RECT 372.120000 412.180000 373.320000 412.660000 ;
        RECT 372.120000 384.980000 373.320000 385.460000 ;
        RECT 372.120000 379.540000 373.320000 380.020000 ;
        RECT 372.120000 390.420000 373.320000 390.900000 ;
        RECT 372.120000 406.740000 373.320000 407.220000 ;
        RECT 372.120000 395.860000 373.320000 396.340000 ;
        RECT 372.120000 401.300000 373.320000 401.780000 ;
        RECT 417.120000 384.980000 418.320000 385.460000 ;
        RECT 417.120000 379.540000 418.320000 380.020000 ;
        RECT 417.120000 390.420000 418.320000 390.900000 ;
        RECT 417.120000 395.860000 418.320000 396.340000 ;
        RECT 417.120000 401.300000 418.320000 401.780000 ;
        RECT 417.120000 406.740000 418.320000 407.220000 ;
        RECT 372.120000 428.500000 373.320000 428.980000 ;
        RECT 372.120000 423.060000 373.320000 423.540000 ;
        RECT 372.120000 417.620000 373.320000 418.100000 ;
        RECT 372.120000 439.380000 373.320000 439.860000 ;
        RECT 372.120000 433.940000 373.320000 434.420000 ;
        RECT 372.120000 444.820000 373.320000 445.300000 ;
        RECT 417.120000 428.500000 418.320000 428.980000 ;
        RECT 417.120000 423.060000 418.320000 423.540000 ;
        RECT 417.120000 417.620000 418.320000 418.100000 ;
        RECT 417.120000 439.380000 418.320000 439.860000 ;
        RECT 417.120000 433.940000 418.320000 434.420000 ;
        RECT 417.120000 444.820000 418.320000 445.300000 ;
        RECT 462.120000 330.580000 463.320000 331.060000 ;
        RECT 462.120000 303.380000 463.320000 303.860000 ;
        RECT 462.120000 308.820000 463.320000 309.300000 ;
        RECT 462.120000 314.260000 463.320000 314.740000 ;
        RECT 462.120000 319.700000 463.320000 320.180000 ;
        RECT 462.120000 325.140000 463.320000 325.620000 ;
        RECT 462.120000 336.020000 463.320000 336.500000 ;
        RECT 462.120000 374.100000 463.320000 374.580000 ;
        RECT 462.120000 368.660000 463.320000 369.140000 ;
        RECT 462.120000 363.220000 463.320000 363.700000 ;
        RECT 462.120000 357.780000 463.320000 358.260000 ;
        RECT 462.120000 341.460000 463.320000 341.940000 ;
        RECT 462.120000 346.900000 463.320000 347.380000 ;
        RECT 462.120000 352.340000 463.320000 352.820000 ;
        RECT 507.120000 303.380000 508.320000 303.860000 ;
        RECT 507.120000 308.820000 508.320000 309.300000 ;
        RECT 507.120000 314.260000 508.320000 314.740000 ;
        RECT 507.120000 319.700000 508.320000 320.180000 ;
        RECT 507.120000 325.140000 508.320000 325.620000 ;
        RECT 507.120000 330.580000 508.320000 331.060000 ;
        RECT 507.120000 336.020000 508.320000 336.500000 ;
        RECT 543.400000 314.260000 544.600000 314.740000 ;
        RECT 543.400000 308.820000 544.600000 309.300000 ;
        RECT 543.400000 303.380000 544.600000 303.860000 ;
        RECT 543.400000 336.020000 544.600000 336.500000 ;
        RECT 543.400000 330.580000 544.600000 331.060000 ;
        RECT 543.400000 325.140000 544.600000 325.620000 ;
        RECT 543.400000 319.700000 544.600000 320.180000 ;
        RECT 507.120000 341.460000 508.320000 341.940000 ;
        RECT 507.120000 346.900000 508.320000 347.380000 ;
        RECT 507.120000 352.340000 508.320000 352.820000 ;
        RECT 507.120000 374.100000 508.320000 374.580000 ;
        RECT 507.120000 368.660000 508.320000 369.140000 ;
        RECT 507.120000 363.220000 508.320000 363.700000 ;
        RECT 507.120000 357.780000 508.320000 358.260000 ;
        RECT 543.400000 352.340000 544.600000 352.820000 ;
        RECT 543.400000 346.900000 544.600000 347.380000 ;
        RECT 543.400000 341.460000 544.600000 341.940000 ;
        RECT 543.400000 374.100000 544.600000 374.580000 ;
        RECT 543.400000 368.660000 544.600000 369.140000 ;
        RECT 543.400000 363.220000 544.600000 363.700000 ;
        RECT 543.400000 357.780000 544.600000 358.260000 ;
        RECT 462.120000 412.180000 463.320000 412.660000 ;
        RECT 462.120000 401.300000 463.320000 401.780000 ;
        RECT 462.120000 395.860000 463.320000 396.340000 ;
        RECT 462.120000 390.420000 463.320000 390.900000 ;
        RECT 462.120000 384.980000 463.320000 385.460000 ;
        RECT 462.120000 379.540000 463.320000 380.020000 ;
        RECT 462.120000 406.740000 463.320000 407.220000 ;
        RECT 462.120000 444.820000 463.320000 445.300000 ;
        RECT 462.120000 439.380000 463.320000 439.860000 ;
        RECT 462.120000 433.940000 463.320000 434.420000 ;
        RECT 462.120000 417.620000 463.320000 418.100000 ;
        RECT 462.120000 423.060000 463.320000 423.540000 ;
        RECT 462.120000 428.500000 463.320000 428.980000 ;
        RECT 543.400000 412.180000 544.600000 412.660000 ;
        RECT 507.120000 412.180000 508.320000 412.660000 ;
        RECT 507.120000 390.420000 508.320000 390.900000 ;
        RECT 507.120000 384.980000 508.320000 385.460000 ;
        RECT 507.120000 379.540000 508.320000 380.020000 ;
        RECT 507.120000 401.300000 508.320000 401.780000 ;
        RECT 507.120000 395.860000 508.320000 396.340000 ;
        RECT 507.120000 406.740000 508.320000 407.220000 ;
        RECT 543.400000 390.420000 544.600000 390.900000 ;
        RECT 543.400000 384.980000 544.600000 385.460000 ;
        RECT 543.400000 379.540000 544.600000 380.020000 ;
        RECT 543.400000 406.740000 544.600000 407.220000 ;
        RECT 543.400000 401.300000 544.600000 401.780000 ;
        RECT 543.400000 395.860000 544.600000 396.340000 ;
        RECT 507.120000 417.620000 508.320000 418.100000 ;
        RECT 507.120000 423.060000 508.320000 423.540000 ;
        RECT 507.120000 428.500000 508.320000 428.980000 ;
        RECT 507.120000 444.820000 508.320000 445.300000 ;
        RECT 507.120000 439.380000 508.320000 439.860000 ;
        RECT 507.120000 433.940000 508.320000 434.420000 ;
        RECT 543.400000 428.500000 544.600000 428.980000 ;
        RECT 543.400000 423.060000 544.600000 423.540000 ;
        RECT 543.400000 417.620000 544.600000 418.100000 ;
        RECT 543.400000 444.820000 544.600000 445.300000 ;
        RECT 543.400000 439.380000 544.600000 439.860000 ;
        RECT 543.400000 433.940000 544.600000 434.420000 ;
        RECT 282.120000 461.140000 283.320000 461.620000 ;
        RECT 282.120000 450.260000 283.320000 450.740000 ;
        RECT 282.120000 455.700000 283.320000 456.180000 ;
        RECT 282.120000 466.580000 283.320000 467.060000 ;
        RECT 282.120000 477.460000 283.320000 477.940000 ;
        RECT 282.120000 472.020000 283.320000 472.500000 ;
        RECT 282.120000 482.900000 283.320000 483.380000 ;
        RECT 327.120000 461.140000 328.320000 461.620000 ;
        RECT 327.120000 450.260000 328.320000 450.740000 ;
        RECT 327.120000 455.700000 328.320000 456.180000 ;
        RECT 327.120000 466.580000 328.320000 467.060000 ;
        RECT 327.120000 472.020000 328.320000 472.500000 ;
        RECT 327.120000 477.460000 328.320000 477.940000 ;
        RECT 327.120000 482.900000 328.320000 483.380000 ;
        RECT 282.120000 504.660000 283.320000 505.140000 ;
        RECT 282.120000 499.220000 283.320000 499.700000 ;
        RECT 282.120000 493.780000 283.320000 494.260000 ;
        RECT 282.120000 488.340000 283.320000 488.820000 ;
        RECT 282.120000 510.100000 283.320000 510.580000 ;
        RECT 282.120000 515.540000 283.320000 516.020000 ;
        RECT 282.120000 520.980000 283.320000 521.460000 ;
        RECT 327.120000 504.660000 328.320000 505.140000 ;
        RECT 327.120000 499.220000 328.320000 499.700000 ;
        RECT 327.120000 493.780000 328.320000 494.260000 ;
        RECT 327.120000 488.340000 328.320000 488.820000 ;
        RECT 327.120000 510.100000 328.320000 510.580000 ;
        RECT 327.120000 515.540000 328.320000 516.020000 ;
        RECT 327.120000 520.980000 328.320000 521.460000 ;
        RECT 372.120000 450.260000 373.320000 450.740000 ;
        RECT 372.120000 455.700000 373.320000 456.180000 ;
        RECT 372.120000 461.140000 373.320000 461.620000 ;
        RECT 372.120000 466.580000 373.320000 467.060000 ;
        RECT 372.120000 477.460000 373.320000 477.940000 ;
        RECT 372.120000 472.020000 373.320000 472.500000 ;
        RECT 372.120000 482.900000 373.320000 483.380000 ;
        RECT 417.120000 450.260000 418.320000 450.740000 ;
        RECT 417.120000 455.700000 418.320000 456.180000 ;
        RECT 417.120000 461.140000 418.320000 461.620000 ;
        RECT 417.120000 466.580000 418.320000 467.060000 ;
        RECT 417.120000 472.020000 418.320000 472.500000 ;
        RECT 417.120000 477.460000 418.320000 477.940000 ;
        RECT 417.120000 482.900000 418.320000 483.380000 ;
        RECT 372.120000 504.660000 373.320000 505.140000 ;
        RECT 372.120000 499.220000 373.320000 499.700000 ;
        RECT 372.120000 493.780000 373.320000 494.260000 ;
        RECT 372.120000 488.340000 373.320000 488.820000 ;
        RECT 372.120000 510.100000 373.320000 510.580000 ;
        RECT 372.120000 515.540000 373.320000 516.020000 ;
        RECT 372.120000 520.980000 373.320000 521.460000 ;
        RECT 417.120000 504.660000 418.320000 505.140000 ;
        RECT 417.120000 499.220000 418.320000 499.700000 ;
        RECT 417.120000 493.780000 418.320000 494.260000 ;
        RECT 417.120000 488.340000 418.320000 488.820000 ;
        RECT 417.120000 510.100000 418.320000 510.580000 ;
        RECT 417.120000 515.540000 418.320000 516.020000 ;
        RECT 417.120000 520.980000 418.320000 521.460000 ;
        RECT 282.120000 531.860000 283.320000 532.340000 ;
        RECT 282.120000 526.420000 283.320000 526.900000 ;
        RECT 282.120000 537.300000 283.320000 537.780000 ;
        RECT 282.120000 542.740000 283.320000 543.220000 ;
        RECT 282.120000 548.180000 283.320000 548.660000 ;
        RECT 282.120000 553.620000 283.320000 554.100000 ;
        RECT 282.120000 559.060000 283.320000 559.540000 ;
        RECT 327.120000 531.860000 328.320000 532.340000 ;
        RECT 327.120000 526.420000 328.320000 526.900000 ;
        RECT 327.120000 537.300000 328.320000 537.780000 ;
        RECT 327.120000 542.740000 328.320000 543.220000 ;
        RECT 327.120000 548.180000 328.320000 548.660000 ;
        RECT 327.120000 553.620000 328.320000 554.100000 ;
        RECT 327.120000 559.060000 328.320000 559.540000 ;
        RECT 282.120000 580.820000 283.320000 581.300000 ;
        RECT 282.120000 575.380000 283.320000 575.860000 ;
        RECT 282.120000 569.940000 283.320000 570.420000 ;
        RECT 282.120000 564.500000 283.320000 564.980000 ;
        RECT 282.120000 586.260000 283.320000 586.740000 ;
        RECT 327.120000 580.820000 328.320000 581.300000 ;
        RECT 327.120000 575.380000 328.320000 575.860000 ;
        RECT 327.120000 569.940000 328.320000 570.420000 ;
        RECT 327.120000 564.500000 328.320000 564.980000 ;
        RECT 327.120000 586.260000 328.320000 586.740000 ;
        RECT 372.120000 531.860000 373.320000 532.340000 ;
        RECT 372.120000 526.420000 373.320000 526.900000 ;
        RECT 372.120000 537.300000 373.320000 537.780000 ;
        RECT 372.120000 542.740000 373.320000 543.220000 ;
        RECT 372.120000 548.180000 373.320000 548.660000 ;
        RECT 372.120000 553.620000 373.320000 554.100000 ;
        RECT 372.120000 559.060000 373.320000 559.540000 ;
        RECT 417.120000 531.860000 418.320000 532.340000 ;
        RECT 417.120000 526.420000 418.320000 526.900000 ;
        RECT 417.120000 537.300000 418.320000 537.780000 ;
        RECT 417.120000 542.740000 418.320000 543.220000 ;
        RECT 417.120000 548.180000 418.320000 548.660000 ;
        RECT 417.120000 553.620000 418.320000 554.100000 ;
        RECT 417.120000 559.060000 418.320000 559.540000 ;
        RECT 372.120000 580.820000 373.320000 581.300000 ;
        RECT 372.120000 575.380000 373.320000 575.860000 ;
        RECT 372.120000 569.940000 373.320000 570.420000 ;
        RECT 372.120000 564.500000 373.320000 564.980000 ;
        RECT 372.120000 586.260000 373.320000 586.740000 ;
        RECT 417.120000 580.820000 418.320000 581.300000 ;
        RECT 417.120000 575.380000 418.320000 575.860000 ;
        RECT 417.120000 569.940000 418.320000 570.420000 ;
        RECT 417.120000 564.500000 418.320000 564.980000 ;
        RECT 417.120000 586.260000 418.320000 586.740000 ;
        RECT 462.120000 472.020000 463.320000 472.500000 ;
        RECT 462.120000 450.260000 463.320000 450.740000 ;
        RECT 462.120000 455.700000 463.320000 456.180000 ;
        RECT 462.120000 461.140000 463.320000 461.620000 ;
        RECT 462.120000 466.580000 463.320000 467.060000 ;
        RECT 462.120000 477.460000 463.320000 477.940000 ;
        RECT 462.120000 482.900000 463.320000 483.380000 ;
        RECT 462.120000 520.980000 463.320000 521.460000 ;
        RECT 462.120000 515.540000 463.320000 516.020000 ;
        RECT 462.120000 510.100000 463.320000 510.580000 ;
        RECT 462.120000 504.660000 463.320000 505.140000 ;
        RECT 462.120000 488.340000 463.320000 488.820000 ;
        RECT 462.120000 493.780000 463.320000 494.260000 ;
        RECT 462.120000 499.220000 463.320000 499.700000 ;
        RECT 507.120000 450.260000 508.320000 450.740000 ;
        RECT 507.120000 455.700000 508.320000 456.180000 ;
        RECT 507.120000 461.140000 508.320000 461.620000 ;
        RECT 507.120000 466.580000 508.320000 467.060000 ;
        RECT 507.120000 472.020000 508.320000 472.500000 ;
        RECT 507.120000 477.460000 508.320000 477.940000 ;
        RECT 507.120000 482.900000 508.320000 483.380000 ;
        RECT 543.400000 466.580000 544.600000 467.060000 ;
        RECT 543.400000 461.140000 544.600000 461.620000 ;
        RECT 543.400000 455.700000 544.600000 456.180000 ;
        RECT 543.400000 450.260000 544.600000 450.740000 ;
        RECT 543.400000 482.900000 544.600000 483.380000 ;
        RECT 543.400000 477.460000 544.600000 477.940000 ;
        RECT 543.400000 472.020000 544.600000 472.500000 ;
        RECT 507.120000 504.660000 508.320000 505.140000 ;
        RECT 507.120000 488.340000 508.320000 488.820000 ;
        RECT 507.120000 493.780000 508.320000 494.260000 ;
        RECT 507.120000 499.220000 508.320000 499.700000 ;
        RECT 507.120000 520.980000 508.320000 521.460000 ;
        RECT 507.120000 515.540000 508.320000 516.020000 ;
        RECT 507.120000 510.100000 508.320000 510.580000 ;
        RECT 543.400000 504.660000 544.600000 505.140000 ;
        RECT 543.400000 499.220000 544.600000 499.700000 ;
        RECT 543.400000 493.780000 544.600000 494.260000 ;
        RECT 543.400000 488.340000 544.600000 488.820000 ;
        RECT 543.400000 520.980000 544.600000 521.460000 ;
        RECT 543.400000 515.540000 544.600000 516.020000 ;
        RECT 543.400000 510.100000 544.600000 510.580000 ;
        RECT 462.120000 542.740000 463.320000 543.220000 ;
        RECT 462.120000 537.300000 463.320000 537.780000 ;
        RECT 462.120000 531.860000 463.320000 532.340000 ;
        RECT 462.120000 526.420000 463.320000 526.900000 ;
        RECT 462.120000 548.180000 463.320000 548.660000 ;
        RECT 462.120000 553.620000 463.320000 554.100000 ;
        RECT 462.120000 559.060000 463.320000 559.540000 ;
        RECT 462.120000 586.260000 463.320000 586.740000 ;
        RECT 462.120000 580.820000 463.320000 581.300000 ;
        RECT 462.120000 564.500000 463.320000 564.980000 ;
        RECT 462.120000 569.940000 463.320000 570.420000 ;
        RECT 462.120000 575.380000 463.320000 575.860000 ;
        RECT 507.120000 542.740000 508.320000 543.220000 ;
        RECT 507.120000 537.300000 508.320000 537.780000 ;
        RECT 507.120000 531.860000 508.320000 532.340000 ;
        RECT 507.120000 526.420000 508.320000 526.900000 ;
        RECT 507.120000 548.180000 508.320000 548.660000 ;
        RECT 507.120000 553.620000 508.320000 554.100000 ;
        RECT 507.120000 559.060000 508.320000 559.540000 ;
        RECT 543.400000 542.740000 544.600000 543.220000 ;
        RECT 543.400000 537.300000 544.600000 537.780000 ;
        RECT 543.400000 531.860000 544.600000 532.340000 ;
        RECT 543.400000 526.420000 544.600000 526.900000 ;
        RECT 543.400000 559.060000 544.600000 559.540000 ;
        RECT 543.400000 553.620000 544.600000 554.100000 ;
        RECT 543.400000 548.180000 544.600000 548.660000 ;
        RECT 507.120000 580.820000 508.320000 581.300000 ;
        RECT 507.120000 575.380000 508.320000 575.860000 ;
        RECT 507.120000 564.500000 508.320000 564.980000 ;
        RECT 507.120000 569.940000 508.320000 570.420000 ;
        RECT 507.120000 586.260000 508.320000 586.740000 ;
        RECT 543.400000 580.820000 544.600000 581.300000 ;
        RECT 543.400000 575.380000 544.600000 575.860000 ;
        RECT 543.400000 569.940000 544.600000 570.420000 ;
        RECT 543.400000 564.500000 544.600000 564.980000 ;
        RECT 543.400000 586.260000 544.600000 586.740000 ;
      LAYER met4 ;
        RECT 507.120000 5.430000 508.320000 593.990000 ;
        RECT 462.120000 5.430000 463.320000 593.990000 ;
        RECT 417.120000 5.430000 418.320000 593.990000 ;
        RECT 372.120000 5.430000 373.320000 593.990000 ;
        RECT 327.120000 5.430000 328.320000 593.990000 ;
        RECT 282.120000 5.430000 283.320000 593.990000 ;
        RECT 237.120000 5.430000 238.320000 593.990000 ;
        RECT 192.120000 5.430000 193.320000 593.990000 ;
        RECT 147.120000 5.430000 148.320000 593.990000 ;
        RECT 102.120000 5.430000 103.320000 593.990000 ;
        RECT 57.120000 5.430000 58.320000 593.990000 ;
        RECT 12.120000 5.430000 13.320000 593.990000 ;
        RECT 543.400000 0.000000 544.600000 599.760000 ;
        RECT 5.560000 0.000000 6.760000 599.760000 ;
    END
# end of P/G power stripe data as pin

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 548.960000 594.990000 550.160000 596.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 594.990000 1.200000 596.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 548.960000 3.230000 550.160000 4.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 3.230000 1.200000 4.430000 ;
    END
    PORT
      LAYER met4 ;
        RECT 545.600000 598.560000 546.800000 599.760000 ;
    END
    PORT
      LAYER met4 ;
        RECT 545.600000 0.000000 546.800000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 3.360000 598.560000 4.560000 599.760000 ;
    END
    PORT
      LAYER met4 ;
        RECT 3.360000 0.000000 4.560000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 3.230000 550.160000 4.430000 ;
        RECT 0.000000 594.990000 550.160000 596.190000 ;
        RECT 3.360000 17.780000 4.560000 18.260000 ;
        RECT 9.955000 17.780000 11.320000 18.260000 ;
        RECT 3.360000 12.340000 4.560000 12.820000 ;
        RECT 9.955000 12.340000 11.320000 12.820000 ;
        RECT 3.360000 23.220000 4.560000 23.700000 ;
        RECT 9.955000 23.220000 11.320000 23.700000 ;
        RECT 3.360000 34.100000 4.560000 34.580000 ;
        RECT 9.955000 34.100000 11.320000 34.580000 ;
        RECT 3.360000 28.660000 4.560000 29.140000 ;
        RECT 9.955000 28.660000 11.320000 29.140000 ;
        RECT 3.360000 55.860000 4.560000 56.340000 ;
        RECT 9.955000 55.860000 11.320000 56.340000 ;
        RECT 3.360000 44.980000 4.560000 45.460000 ;
        RECT 9.955000 44.980000 11.320000 45.460000 ;
        RECT 3.360000 39.540000 4.560000 40.020000 ;
        RECT 9.955000 39.540000 11.320000 40.020000 ;
        RECT 3.360000 50.420000 4.560000 50.900000 ;
        RECT 9.955000 50.420000 11.320000 50.900000 ;
        RECT 3.360000 61.300000 4.560000 61.780000 ;
        RECT 9.955000 61.300000 11.320000 61.780000 ;
        RECT 3.360000 72.180000 4.560000 72.660000 ;
        RECT 3.360000 66.740000 4.560000 67.220000 ;
        RECT 9.955000 66.740000 11.320000 67.220000 ;
        RECT 9.955000 72.180000 11.320000 72.660000 ;
        RECT 55.120000 12.340000 56.320000 12.820000 ;
        RECT 55.120000 17.780000 56.320000 18.260000 ;
        RECT 55.120000 34.100000 56.320000 34.580000 ;
        RECT 55.120000 23.220000 56.320000 23.700000 ;
        RECT 55.120000 28.660000 56.320000 29.140000 ;
        RECT 100.120000 12.340000 101.320000 12.820000 ;
        RECT 100.120000 17.780000 101.320000 18.260000 ;
        RECT 100.120000 34.100000 101.320000 34.580000 ;
        RECT 100.120000 23.220000 101.320000 23.700000 ;
        RECT 100.120000 28.660000 101.320000 29.140000 ;
        RECT 55.120000 55.860000 56.320000 56.340000 ;
        RECT 55.120000 39.540000 56.320000 40.020000 ;
        RECT 55.120000 44.980000 56.320000 45.460000 ;
        RECT 55.120000 50.420000 56.320000 50.900000 ;
        RECT 55.120000 72.180000 56.320000 72.660000 ;
        RECT 55.120000 66.740000 56.320000 67.220000 ;
        RECT 55.120000 61.300000 56.320000 61.780000 ;
        RECT 100.120000 55.860000 101.320000 56.340000 ;
        RECT 100.120000 39.540000 101.320000 40.020000 ;
        RECT 100.120000 44.980000 101.320000 45.460000 ;
        RECT 100.120000 50.420000 101.320000 50.900000 ;
        RECT 100.120000 72.180000 101.320000 72.660000 ;
        RECT 100.120000 66.740000 101.320000 67.220000 ;
        RECT 100.120000 61.300000 101.320000 61.780000 ;
        RECT 3.360000 83.060000 4.560000 83.540000 ;
        RECT 9.955000 83.060000 11.320000 83.540000 ;
        RECT 3.360000 77.620000 4.560000 78.100000 ;
        RECT 9.955000 77.620000 11.320000 78.100000 ;
        RECT 3.360000 88.500000 4.560000 88.980000 ;
        RECT 9.955000 88.500000 11.320000 88.980000 ;
        RECT 3.360000 99.380000 4.560000 99.860000 ;
        RECT 9.955000 99.380000 11.320000 99.860000 ;
        RECT 3.360000 93.940000 4.560000 94.420000 ;
        RECT 9.955000 93.940000 11.320000 94.420000 ;
        RECT 3.360000 110.260000 4.560000 110.740000 ;
        RECT 9.955000 110.260000 11.320000 110.740000 ;
        RECT 3.360000 104.820000 4.560000 105.300000 ;
        RECT 9.955000 104.820000 11.320000 105.300000 ;
        RECT 3.360000 121.140000 4.560000 121.620000 ;
        RECT 3.360000 115.700000 4.560000 116.180000 ;
        RECT 9.955000 115.700000 11.320000 116.180000 ;
        RECT 9.955000 121.140000 11.320000 121.620000 ;
        RECT 3.360000 126.580000 4.560000 127.060000 ;
        RECT 9.955000 126.580000 11.320000 127.060000 ;
        RECT 3.360000 137.460000 4.560000 137.940000 ;
        RECT 9.955000 137.460000 11.320000 137.940000 ;
        RECT 3.360000 132.020000 4.560000 132.500000 ;
        RECT 9.955000 132.020000 11.320000 132.500000 ;
        RECT 3.360000 148.340000 4.560000 148.820000 ;
        RECT 9.955000 148.340000 11.320000 148.820000 ;
        RECT 3.360000 142.900000 4.560000 143.380000 ;
        RECT 9.955000 142.900000 11.320000 143.380000 ;
        RECT 55.120000 77.620000 56.320000 78.100000 ;
        RECT 55.120000 83.060000 56.320000 83.540000 ;
        RECT 55.120000 88.500000 56.320000 88.980000 ;
        RECT 55.120000 110.260000 56.320000 110.740000 ;
        RECT 55.120000 104.820000 56.320000 105.300000 ;
        RECT 55.120000 99.380000 56.320000 99.860000 ;
        RECT 55.120000 93.940000 56.320000 94.420000 ;
        RECT 100.120000 77.620000 101.320000 78.100000 ;
        RECT 100.120000 83.060000 101.320000 83.540000 ;
        RECT 100.120000 88.500000 101.320000 88.980000 ;
        RECT 100.120000 110.260000 101.320000 110.740000 ;
        RECT 100.120000 104.820000 101.320000 105.300000 ;
        RECT 100.120000 99.380000 101.320000 99.860000 ;
        RECT 100.120000 93.940000 101.320000 94.420000 ;
        RECT 55.120000 115.700000 56.320000 116.180000 ;
        RECT 55.120000 121.140000 56.320000 121.620000 ;
        RECT 55.120000 126.580000 56.320000 127.060000 ;
        RECT 55.120000 148.340000 56.320000 148.820000 ;
        RECT 55.120000 142.900000 56.320000 143.380000 ;
        RECT 55.120000 137.460000 56.320000 137.940000 ;
        RECT 55.120000 132.020000 56.320000 132.500000 ;
        RECT 100.120000 115.700000 101.320000 116.180000 ;
        RECT 100.120000 121.140000 101.320000 121.620000 ;
        RECT 100.120000 126.580000 101.320000 127.060000 ;
        RECT 100.120000 148.340000 101.320000 148.820000 ;
        RECT 100.120000 142.900000 101.320000 143.380000 ;
        RECT 100.120000 137.460000 101.320000 137.940000 ;
        RECT 100.120000 132.020000 101.320000 132.500000 ;
        RECT 145.120000 12.340000 146.320000 12.820000 ;
        RECT 145.120000 17.780000 146.320000 18.260000 ;
        RECT 145.120000 34.100000 146.320000 34.580000 ;
        RECT 145.120000 23.220000 146.320000 23.700000 ;
        RECT 145.120000 28.660000 146.320000 29.140000 ;
        RECT 190.120000 12.340000 191.320000 12.820000 ;
        RECT 190.120000 17.780000 191.320000 18.260000 ;
        RECT 190.120000 34.100000 191.320000 34.580000 ;
        RECT 190.120000 23.220000 191.320000 23.700000 ;
        RECT 190.120000 28.660000 191.320000 29.140000 ;
        RECT 145.120000 55.860000 146.320000 56.340000 ;
        RECT 145.120000 39.540000 146.320000 40.020000 ;
        RECT 145.120000 44.980000 146.320000 45.460000 ;
        RECT 145.120000 50.420000 146.320000 50.900000 ;
        RECT 145.120000 72.180000 146.320000 72.660000 ;
        RECT 145.120000 66.740000 146.320000 67.220000 ;
        RECT 145.120000 61.300000 146.320000 61.780000 ;
        RECT 190.120000 55.860000 191.320000 56.340000 ;
        RECT 190.120000 39.540000 191.320000 40.020000 ;
        RECT 190.120000 44.980000 191.320000 45.460000 ;
        RECT 190.120000 50.420000 191.320000 50.900000 ;
        RECT 190.120000 72.180000 191.320000 72.660000 ;
        RECT 190.120000 66.740000 191.320000 67.220000 ;
        RECT 190.120000 61.300000 191.320000 61.780000 ;
        RECT 235.120000 34.100000 236.320000 34.580000 ;
        RECT 235.120000 12.340000 236.320000 12.820000 ;
        RECT 235.120000 17.780000 236.320000 18.260000 ;
        RECT 235.120000 23.220000 236.320000 23.700000 ;
        RECT 235.120000 28.660000 236.320000 29.140000 ;
        RECT 235.120000 72.180000 236.320000 72.660000 ;
        RECT 235.120000 66.740000 236.320000 67.220000 ;
        RECT 235.120000 61.300000 236.320000 61.780000 ;
        RECT 235.120000 39.540000 236.320000 40.020000 ;
        RECT 235.120000 44.980000 236.320000 45.460000 ;
        RECT 235.120000 50.420000 236.320000 50.900000 ;
        RECT 235.120000 55.860000 236.320000 56.340000 ;
        RECT 145.120000 77.620000 146.320000 78.100000 ;
        RECT 145.120000 83.060000 146.320000 83.540000 ;
        RECT 145.120000 88.500000 146.320000 88.980000 ;
        RECT 145.120000 110.260000 146.320000 110.740000 ;
        RECT 145.120000 104.820000 146.320000 105.300000 ;
        RECT 145.120000 99.380000 146.320000 99.860000 ;
        RECT 145.120000 93.940000 146.320000 94.420000 ;
        RECT 190.120000 77.620000 191.320000 78.100000 ;
        RECT 190.120000 83.060000 191.320000 83.540000 ;
        RECT 190.120000 88.500000 191.320000 88.980000 ;
        RECT 190.120000 110.260000 191.320000 110.740000 ;
        RECT 190.120000 104.820000 191.320000 105.300000 ;
        RECT 190.120000 99.380000 191.320000 99.860000 ;
        RECT 190.120000 93.940000 191.320000 94.420000 ;
        RECT 145.120000 115.700000 146.320000 116.180000 ;
        RECT 145.120000 121.140000 146.320000 121.620000 ;
        RECT 145.120000 126.580000 146.320000 127.060000 ;
        RECT 145.120000 148.340000 146.320000 148.820000 ;
        RECT 145.120000 142.900000 146.320000 143.380000 ;
        RECT 145.120000 137.460000 146.320000 137.940000 ;
        RECT 145.120000 132.020000 146.320000 132.500000 ;
        RECT 190.120000 115.700000 191.320000 116.180000 ;
        RECT 190.120000 121.140000 191.320000 121.620000 ;
        RECT 190.120000 126.580000 191.320000 127.060000 ;
        RECT 190.120000 148.340000 191.320000 148.820000 ;
        RECT 190.120000 142.900000 191.320000 143.380000 ;
        RECT 190.120000 137.460000 191.320000 137.940000 ;
        RECT 190.120000 132.020000 191.320000 132.500000 ;
        RECT 235.120000 110.260000 236.320000 110.740000 ;
        RECT 235.120000 104.820000 236.320000 105.300000 ;
        RECT 235.120000 99.380000 236.320000 99.860000 ;
        RECT 235.120000 77.620000 236.320000 78.100000 ;
        RECT 235.120000 83.060000 236.320000 83.540000 ;
        RECT 235.120000 88.500000 236.320000 88.980000 ;
        RECT 235.120000 93.940000 236.320000 94.420000 ;
        RECT 235.120000 148.340000 236.320000 148.820000 ;
        RECT 235.120000 142.900000 236.320000 143.380000 ;
        RECT 235.120000 137.460000 236.320000 137.940000 ;
        RECT 235.120000 132.020000 236.320000 132.500000 ;
        RECT 235.120000 115.700000 236.320000 116.180000 ;
        RECT 235.120000 121.140000 236.320000 121.620000 ;
        RECT 235.120000 126.580000 236.320000 127.060000 ;
        RECT 3.360000 224.500000 4.560000 224.980000 ;
        RECT 9.955000 224.500000 11.320000 224.980000 ;
        RECT 100.120000 224.500000 101.320000 224.980000 ;
        RECT 55.120000 224.500000 56.320000 224.980000 ;
        RECT 3.360000 159.220000 4.560000 159.700000 ;
        RECT 9.955000 159.220000 11.320000 159.700000 ;
        RECT 3.360000 153.780000 4.560000 154.260000 ;
        RECT 9.955000 153.780000 11.320000 154.260000 ;
        RECT 3.360000 164.660000 4.560000 165.140000 ;
        RECT 9.955000 164.660000 11.320000 165.140000 ;
        RECT 3.360000 175.540000 4.560000 176.020000 ;
        RECT 9.955000 175.540000 11.320000 176.020000 ;
        RECT 3.360000 170.100000 4.560000 170.580000 ;
        RECT 9.955000 170.100000 11.320000 170.580000 ;
        RECT 3.360000 186.420000 4.560000 186.900000 ;
        RECT 9.955000 186.420000 11.320000 186.900000 ;
        RECT 3.360000 180.980000 4.560000 181.460000 ;
        RECT 9.955000 180.980000 11.320000 181.460000 ;
        RECT 3.360000 191.860000 4.560000 192.340000 ;
        RECT 9.955000 191.860000 11.320000 192.340000 ;
        RECT 3.360000 202.740000 4.560000 203.220000 ;
        RECT 9.955000 202.740000 11.320000 203.220000 ;
        RECT 3.360000 197.300000 4.560000 197.780000 ;
        RECT 9.955000 197.300000 11.320000 197.780000 ;
        RECT 3.360000 213.620000 4.560000 214.100000 ;
        RECT 9.955000 213.620000 11.320000 214.100000 ;
        RECT 3.360000 208.180000 4.560000 208.660000 ;
        RECT 9.955000 208.180000 11.320000 208.660000 ;
        RECT 3.360000 219.060000 4.560000 219.540000 ;
        RECT 9.955000 219.060000 11.320000 219.540000 ;
        RECT 55.120000 153.780000 56.320000 154.260000 ;
        RECT 55.120000 159.220000 56.320000 159.700000 ;
        RECT 55.120000 164.660000 56.320000 165.140000 ;
        RECT 55.120000 186.420000 56.320000 186.900000 ;
        RECT 55.120000 180.980000 56.320000 181.460000 ;
        RECT 55.120000 175.540000 56.320000 176.020000 ;
        RECT 55.120000 170.100000 56.320000 170.580000 ;
        RECT 100.120000 153.780000 101.320000 154.260000 ;
        RECT 100.120000 159.220000 101.320000 159.700000 ;
        RECT 100.120000 164.660000 101.320000 165.140000 ;
        RECT 100.120000 186.420000 101.320000 186.900000 ;
        RECT 100.120000 180.980000 101.320000 181.460000 ;
        RECT 100.120000 175.540000 101.320000 176.020000 ;
        RECT 100.120000 170.100000 101.320000 170.580000 ;
        RECT 55.120000 191.860000 56.320000 192.340000 ;
        RECT 55.120000 197.300000 56.320000 197.780000 ;
        RECT 55.120000 202.740000 56.320000 203.220000 ;
        RECT 55.120000 219.060000 56.320000 219.540000 ;
        RECT 55.120000 213.620000 56.320000 214.100000 ;
        RECT 55.120000 208.180000 56.320000 208.660000 ;
        RECT 100.120000 191.860000 101.320000 192.340000 ;
        RECT 100.120000 197.300000 101.320000 197.780000 ;
        RECT 100.120000 202.740000 101.320000 203.220000 ;
        RECT 100.120000 219.060000 101.320000 219.540000 ;
        RECT 100.120000 213.620000 101.320000 214.100000 ;
        RECT 100.120000 208.180000 101.320000 208.660000 ;
        RECT 3.360000 229.940000 4.560000 230.420000 ;
        RECT 9.955000 229.940000 11.320000 230.420000 ;
        RECT 3.360000 240.820000 4.560000 241.300000 ;
        RECT 3.360000 235.380000 4.560000 235.860000 ;
        RECT 9.955000 235.380000 11.320000 235.860000 ;
        RECT 9.955000 240.820000 11.320000 241.300000 ;
        RECT 3.360000 251.700000 4.560000 252.180000 ;
        RECT 9.955000 251.700000 11.320000 252.180000 ;
        RECT 3.360000 246.260000 4.560000 246.740000 ;
        RECT 9.955000 246.260000 11.320000 246.740000 ;
        RECT 3.360000 257.140000 4.560000 257.620000 ;
        RECT 9.955000 257.140000 11.320000 257.620000 ;
        RECT 3.360000 268.020000 4.560000 268.500000 ;
        RECT 9.955000 268.020000 11.320000 268.500000 ;
        RECT 3.360000 262.580000 4.560000 263.060000 ;
        RECT 9.955000 262.580000 11.320000 263.060000 ;
        RECT 3.360000 278.900000 4.560000 279.380000 ;
        RECT 9.955000 278.900000 11.320000 279.380000 ;
        RECT 3.360000 273.460000 4.560000 273.940000 ;
        RECT 9.955000 273.460000 11.320000 273.940000 ;
        RECT 3.360000 289.780000 4.560000 290.260000 ;
        RECT 3.360000 284.340000 4.560000 284.820000 ;
        RECT 9.955000 284.340000 11.320000 284.820000 ;
        RECT 9.955000 289.780000 11.320000 290.260000 ;
        RECT 3.360000 295.220000 4.560000 295.700000 ;
        RECT 9.955000 295.220000 11.320000 295.700000 ;
        RECT 55.120000 229.940000 56.320000 230.420000 ;
        RECT 55.120000 235.380000 56.320000 235.860000 ;
        RECT 55.120000 240.820000 56.320000 241.300000 ;
        RECT 55.120000 257.140000 56.320000 257.620000 ;
        RECT 55.120000 251.700000 56.320000 252.180000 ;
        RECT 55.120000 246.260000 56.320000 246.740000 ;
        RECT 100.120000 229.940000 101.320000 230.420000 ;
        RECT 100.120000 235.380000 101.320000 235.860000 ;
        RECT 100.120000 240.820000 101.320000 241.300000 ;
        RECT 100.120000 257.140000 101.320000 257.620000 ;
        RECT 100.120000 251.700000 101.320000 252.180000 ;
        RECT 100.120000 246.260000 101.320000 246.740000 ;
        RECT 55.120000 278.900000 56.320000 279.380000 ;
        RECT 55.120000 262.580000 56.320000 263.060000 ;
        RECT 55.120000 268.020000 56.320000 268.500000 ;
        RECT 55.120000 273.460000 56.320000 273.940000 ;
        RECT 55.120000 295.220000 56.320000 295.700000 ;
        RECT 55.120000 289.780000 56.320000 290.260000 ;
        RECT 55.120000 284.340000 56.320000 284.820000 ;
        RECT 100.120000 278.900000 101.320000 279.380000 ;
        RECT 100.120000 262.580000 101.320000 263.060000 ;
        RECT 100.120000 268.020000 101.320000 268.500000 ;
        RECT 100.120000 273.460000 101.320000 273.940000 ;
        RECT 100.120000 295.220000 101.320000 295.700000 ;
        RECT 100.120000 289.780000 101.320000 290.260000 ;
        RECT 100.120000 284.340000 101.320000 284.820000 ;
        RECT 190.120000 224.500000 191.320000 224.980000 ;
        RECT 145.120000 224.500000 146.320000 224.980000 ;
        RECT 235.120000 224.500000 236.320000 224.980000 ;
        RECT 145.120000 153.780000 146.320000 154.260000 ;
        RECT 145.120000 159.220000 146.320000 159.700000 ;
        RECT 145.120000 164.660000 146.320000 165.140000 ;
        RECT 145.120000 186.420000 146.320000 186.900000 ;
        RECT 145.120000 180.980000 146.320000 181.460000 ;
        RECT 145.120000 175.540000 146.320000 176.020000 ;
        RECT 145.120000 170.100000 146.320000 170.580000 ;
        RECT 190.120000 153.780000 191.320000 154.260000 ;
        RECT 190.120000 159.220000 191.320000 159.700000 ;
        RECT 190.120000 164.660000 191.320000 165.140000 ;
        RECT 190.120000 186.420000 191.320000 186.900000 ;
        RECT 190.120000 180.980000 191.320000 181.460000 ;
        RECT 190.120000 175.540000 191.320000 176.020000 ;
        RECT 190.120000 170.100000 191.320000 170.580000 ;
        RECT 145.120000 191.860000 146.320000 192.340000 ;
        RECT 145.120000 197.300000 146.320000 197.780000 ;
        RECT 145.120000 202.740000 146.320000 203.220000 ;
        RECT 145.120000 219.060000 146.320000 219.540000 ;
        RECT 145.120000 213.620000 146.320000 214.100000 ;
        RECT 145.120000 208.180000 146.320000 208.660000 ;
        RECT 190.120000 191.860000 191.320000 192.340000 ;
        RECT 190.120000 197.300000 191.320000 197.780000 ;
        RECT 190.120000 202.740000 191.320000 203.220000 ;
        RECT 190.120000 219.060000 191.320000 219.540000 ;
        RECT 190.120000 213.620000 191.320000 214.100000 ;
        RECT 190.120000 208.180000 191.320000 208.660000 ;
        RECT 235.120000 186.420000 236.320000 186.900000 ;
        RECT 235.120000 180.980000 236.320000 181.460000 ;
        RECT 235.120000 175.540000 236.320000 176.020000 ;
        RECT 235.120000 170.100000 236.320000 170.580000 ;
        RECT 235.120000 153.780000 236.320000 154.260000 ;
        RECT 235.120000 159.220000 236.320000 159.700000 ;
        RECT 235.120000 164.660000 236.320000 165.140000 ;
        RECT 235.120000 219.060000 236.320000 219.540000 ;
        RECT 235.120000 213.620000 236.320000 214.100000 ;
        RECT 235.120000 208.180000 236.320000 208.660000 ;
        RECT 235.120000 191.860000 236.320000 192.340000 ;
        RECT 235.120000 197.300000 236.320000 197.780000 ;
        RECT 235.120000 202.740000 236.320000 203.220000 ;
        RECT 145.120000 229.940000 146.320000 230.420000 ;
        RECT 145.120000 235.380000 146.320000 235.860000 ;
        RECT 145.120000 240.820000 146.320000 241.300000 ;
        RECT 145.120000 257.140000 146.320000 257.620000 ;
        RECT 145.120000 251.700000 146.320000 252.180000 ;
        RECT 145.120000 246.260000 146.320000 246.740000 ;
        RECT 190.120000 229.940000 191.320000 230.420000 ;
        RECT 190.120000 235.380000 191.320000 235.860000 ;
        RECT 190.120000 240.820000 191.320000 241.300000 ;
        RECT 190.120000 257.140000 191.320000 257.620000 ;
        RECT 190.120000 251.700000 191.320000 252.180000 ;
        RECT 190.120000 246.260000 191.320000 246.740000 ;
        RECT 145.120000 278.900000 146.320000 279.380000 ;
        RECT 145.120000 262.580000 146.320000 263.060000 ;
        RECT 145.120000 268.020000 146.320000 268.500000 ;
        RECT 145.120000 273.460000 146.320000 273.940000 ;
        RECT 145.120000 295.220000 146.320000 295.700000 ;
        RECT 145.120000 289.780000 146.320000 290.260000 ;
        RECT 145.120000 284.340000 146.320000 284.820000 ;
        RECT 190.120000 278.900000 191.320000 279.380000 ;
        RECT 190.120000 262.580000 191.320000 263.060000 ;
        RECT 190.120000 268.020000 191.320000 268.500000 ;
        RECT 190.120000 273.460000 191.320000 273.940000 ;
        RECT 190.120000 295.220000 191.320000 295.700000 ;
        RECT 190.120000 289.780000 191.320000 290.260000 ;
        RECT 190.120000 284.340000 191.320000 284.820000 ;
        RECT 235.120000 257.140000 236.320000 257.620000 ;
        RECT 235.120000 251.700000 236.320000 252.180000 ;
        RECT 235.120000 246.260000 236.320000 246.740000 ;
        RECT 235.120000 229.940000 236.320000 230.420000 ;
        RECT 235.120000 235.380000 236.320000 235.860000 ;
        RECT 235.120000 240.820000 236.320000 241.300000 ;
        RECT 235.120000 295.220000 236.320000 295.700000 ;
        RECT 235.120000 289.780000 236.320000 290.260000 ;
        RECT 235.120000 284.340000 236.320000 284.820000 ;
        RECT 235.120000 278.900000 236.320000 279.380000 ;
        RECT 235.120000 262.580000 236.320000 263.060000 ;
        RECT 235.120000 268.020000 236.320000 268.500000 ;
        RECT 235.120000 273.460000 236.320000 273.940000 ;
        RECT 280.120000 12.340000 281.320000 12.820000 ;
        RECT 280.120000 17.780000 281.320000 18.260000 ;
        RECT 280.120000 34.100000 281.320000 34.580000 ;
        RECT 280.120000 23.220000 281.320000 23.700000 ;
        RECT 280.120000 28.660000 281.320000 29.140000 ;
        RECT 325.120000 12.340000 326.320000 12.820000 ;
        RECT 325.120000 17.780000 326.320000 18.260000 ;
        RECT 325.120000 34.100000 326.320000 34.580000 ;
        RECT 325.120000 23.220000 326.320000 23.700000 ;
        RECT 325.120000 28.660000 326.320000 29.140000 ;
        RECT 280.120000 55.860000 281.320000 56.340000 ;
        RECT 280.120000 39.540000 281.320000 40.020000 ;
        RECT 280.120000 44.980000 281.320000 45.460000 ;
        RECT 280.120000 50.420000 281.320000 50.900000 ;
        RECT 280.120000 72.180000 281.320000 72.660000 ;
        RECT 280.120000 66.740000 281.320000 67.220000 ;
        RECT 280.120000 61.300000 281.320000 61.780000 ;
        RECT 325.120000 55.860000 326.320000 56.340000 ;
        RECT 325.120000 39.540000 326.320000 40.020000 ;
        RECT 325.120000 44.980000 326.320000 45.460000 ;
        RECT 325.120000 50.420000 326.320000 50.900000 ;
        RECT 325.120000 72.180000 326.320000 72.660000 ;
        RECT 325.120000 66.740000 326.320000 67.220000 ;
        RECT 325.120000 61.300000 326.320000 61.780000 ;
        RECT 370.120000 12.340000 371.320000 12.820000 ;
        RECT 370.120000 17.780000 371.320000 18.260000 ;
        RECT 370.120000 34.100000 371.320000 34.580000 ;
        RECT 370.120000 23.220000 371.320000 23.700000 ;
        RECT 370.120000 28.660000 371.320000 29.140000 ;
        RECT 415.120000 12.340000 416.320000 12.820000 ;
        RECT 415.120000 17.780000 416.320000 18.260000 ;
        RECT 415.120000 34.100000 416.320000 34.580000 ;
        RECT 415.120000 23.220000 416.320000 23.700000 ;
        RECT 415.120000 28.660000 416.320000 29.140000 ;
        RECT 370.120000 55.860000 371.320000 56.340000 ;
        RECT 370.120000 39.540000 371.320000 40.020000 ;
        RECT 370.120000 44.980000 371.320000 45.460000 ;
        RECT 370.120000 50.420000 371.320000 50.900000 ;
        RECT 370.120000 72.180000 371.320000 72.660000 ;
        RECT 370.120000 66.740000 371.320000 67.220000 ;
        RECT 370.120000 61.300000 371.320000 61.780000 ;
        RECT 415.120000 55.860000 416.320000 56.340000 ;
        RECT 415.120000 39.540000 416.320000 40.020000 ;
        RECT 415.120000 44.980000 416.320000 45.460000 ;
        RECT 415.120000 50.420000 416.320000 50.900000 ;
        RECT 415.120000 72.180000 416.320000 72.660000 ;
        RECT 415.120000 66.740000 416.320000 67.220000 ;
        RECT 415.120000 61.300000 416.320000 61.780000 ;
        RECT 280.120000 77.620000 281.320000 78.100000 ;
        RECT 280.120000 83.060000 281.320000 83.540000 ;
        RECT 280.120000 88.500000 281.320000 88.980000 ;
        RECT 280.120000 110.260000 281.320000 110.740000 ;
        RECT 280.120000 104.820000 281.320000 105.300000 ;
        RECT 280.120000 99.380000 281.320000 99.860000 ;
        RECT 280.120000 93.940000 281.320000 94.420000 ;
        RECT 325.120000 77.620000 326.320000 78.100000 ;
        RECT 325.120000 83.060000 326.320000 83.540000 ;
        RECT 325.120000 88.500000 326.320000 88.980000 ;
        RECT 325.120000 110.260000 326.320000 110.740000 ;
        RECT 325.120000 104.820000 326.320000 105.300000 ;
        RECT 325.120000 99.380000 326.320000 99.860000 ;
        RECT 325.120000 93.940000 326.320000 94.420000 ;
        RECT 280.120000 115.700000 281.320000 116.180000 ;
        RECT 280.120000 121.140000 281.320000 121.620000 ;
        RECT 280.120000 126.580000 281.320000 127.060000 ;
        RECT 280.120000 148.340000 281.320000 148.820000 ;
        RECT 280.120000 142.900000 281.320000 143.380000 ;
        RECT 280.120000 137.460000 281.320000 137.940000 ;
        RECT 280.120000 132.020000 281.320000 132.500000 ;
        RECT 325.120000 115.700000 326.320000 116.180000 ;
        RECT 325.120000 121.140000 326.320000 121.620000 ;
        RECT 325.120000 126.580000 326.320000 127.060000 ;
        RECT 325.120000 148.340000 326.320000 148.820000 ;
        RECT 325.120000 142.900000 326.320000 143.380000 ;
        RECT 325.120000 137.460000 326.320000 137.940000 ;
        RECT 325.120000 132.020000 326.320000 132.500000 ;
        RECT 370.120000 77.620000 371.320000 78.100000 ;
        RECT 370.120000 83.060000 371.320000 83.540000 ;
        RECT 370.120000 88.500000 371.320000 88.980000 ;
        RECT 370.120000 110.260000 371.320000 110.740000 ;
        RECT 370.120000 104.820000 371.320000 105.300000 ;
        RECT 370.120000 99.380000 371.320000 99.860000 ;
        RECT 370.120000 93.940000 371.320000 94.420000 ;
        RECT 415.120000 77.620000 416.320000 78.100000 ;
        RECT 415.120000 83.060000 416.320000 83.540000 ;
        RECT 415.120000 88.500000 416.320000 88.980000 ;
        RECT 415.120000 110.260000 416.320000 110.740000 ;
        RECT 415.120000 104.820000 416.320000 105.300000 ;
        RECT 415.120000 99.380000 416.320000 99.860000 ;
        RECT 415.120000 93.940000 416.320000 94.420000 ;
        RECT 370.120000 115.700000 371.320000 116.180000 ;
        RECT 370.120000 121.140000 371.320000 121.620000 ;
        RECT 370.120000 126.580000 371.320000 127.060000 ;
        RECT 370.120000 148.340000 371.320000 148.820000 ;
        RECT 370.120000 142.900000 371.320000 143.380000 ;
        RECT 370.120000 137.460000 371.320000 137.940000 ;
        RECT 370.120000 132.020000 371.320000 132.500000 ;
        RECT 415.120000 115.700000 416.320000 116.180000 ;
        RECT 415.120000 121.140000 416.320000 121.620000 ;
        RECT 415.120000 126.580000 416.320000 127.060000 ;
        RECT 415.120000 148.340000 416.320000 148.820000 ;
        RECT 415.120000 142.900000 416.320000 143.380000 ;
        RECT 415.120000 137.460000 416.320000 137.940000 ;
        RECT 415.120000 132.020000 416.320000 132.500000 ;
        RECT 460.120000 34.100000 461.320000 34.580000 ;
        RECT 460.120000 12.340000 461.320000 12.820000 ;
        RECT 460.120000 17.780000 461.320000 18.260000 ;
        RECT 460.120000 23.220000 461.320000 23.700000 ;
        RECT 460.120000 28.660000 461.320000 29.140000 ;
        RECT 460.120000 72.180000 461.320000 72.660000 ;
        RECT 460.120000 66.740000 461.320000 67.220000 ;
        RECT 460.120000 61.300000 461.320000 61.780000 ;
        RECT 460.120000 39.540000 461.320000 40.020000 ;
        RECT 460.120000 44.980000 461.320000 45.460000 ;
        RECT 460.120000 50.420000 461.320000 50.900000 ;
        RECT 460.120000 55.860000 461.320000 56.340000 ;
        RECT 505.120000 17.780000 506.320000 18.260000 ;
        RECT 505.120000 12.340000 506.320000 12.820000 ;
        RECT 505.120000 34.100000 506.320000 34.580000 ;
        RECT 505.120000 23.220000 506.320000 23.700000 ;
        RECT 505.120000 28.660000 506.320000 29.140000 ;
        RECT 545.600000 17.780000 546.800000 18.260000 ;
        RECT 545.600000 12.340000 546.800000 12.820000 ;
        RECT 545.600000 34.100000 546.800000 34.580000 ;
        RECT 545.600000 28.660000 546.800000 29.140000 ;
        RECT 545.600000 23.220000 546.800000 23.700000 ;
        RECT 505.120000 55.860000 506.320000 56.340000 ;
        RECT 505.120000 50.420000 506.320000 50.900000 ;
        RECT 505.120000 44.980000 506.320000 45.460000 ;
        RECT 505.120000 39.540000 506.320000 40.020000 ;
        RECT 505.120000 72.180000 506.320000 72.660000 ;
        RECT 505.120000 66.740000 506.320000 67.220000 ;
        RECT 505.120000 61.300000 506.320000 61.780000 ;
        RECT 545.600000 55.860000 546.800000 56.340000 ;
        RECT 545.600000 50.420000 546.800000 50.900000 ;
        RECT 545.600000 39.540000 546.800000 40.020000 ;
        RECT 545.600000 44.980000 546.800000 45.460000 ;
        RECT 545.600000 72.180000 546.800000 72.660000 ;
        RECT 545.600000 66.740000 546.800000 67.220000 ;
        RECT 545.600000 61.300000 546.800000 61.780000 ;
        RECT 460.120000 110.260000 461.320000 110.740000 ;
        RECT 460.120000 104.820000 461.320000 105.300000 ;
        RECT 460.120000 99.380000 461.320000 99.860000 ;
        RECT 460.120000 77.620000 461.320000 78.100000 ;
        RECT 460.120000 83.060000 461.320000 83.540000 ;
        RECT 460.120000 88.500000 461.320000 88.980000 ;
        RECT 460.120000 93.940000 461.320000 94.420000 ;
        RECT 460.120000 148.340000 461.320000 148.820000 ;
        RECT 460.120000 142.900000 461.320000 143.380000 ;
        RECT 460.120000 137.460000 461.320000 137.940000 ;
        RECT 460.120000 132.020000 461.320000 132.500000 ;
        RECT 460.120000 115.700000 461.320000 116.180000 ;
        RECT 460.120000 121.140000 461.320000 121.620000 ;
        RECT 460.120000 126.580000 461.320000 127.060000 ;
        RECT 505.120000 88.500000 506.320000 88.980000 ;
        RECT 505.120000 83.060000 506.320000 83.540000 ;
        RECT 505.120000 77.620000 506.320000 78.100000 ;
        RECT 505.120000 110.260000 506.320000 110.740000 ;
        RECT 505.120000 104.820000 506.320000 105.300000 ;
        RECT 505.120000 93.940000 506.320000 94.420000 ;
        RECT 505.120000 99.380000 506.320000 99.860000 ;
        RECT 545.600000 88.500000 546.800000 88.980000 ;
        RECT 545.600000 77.620000 546.800000 78.100000 ;
        RECT 545.600000 83.060000 546.800000 83.540000 ;
        RECT 545.600000 110.260000 546.800000 110.740000 ;
        RECT 545.600000 104.820000 546.800000 105.300000 ;
        RECT 545.600000 99.380000 546.800000 99.860000 ;
        RECT 545.600000 93.940000 546.800000 94.420000 ;
        RECT 505.120000 126.580000 506.320000 127.060000 ;
        RECT 505.120000 121.140000 506.320000 121.620000 ;
        RECT 505.120000 115.700000 506.320000 116.180000 ;
        RECT 505.120000 148.340000 506.320000 148.820000 ;
        RECT 505.120000 142.900000 506.320000 143.380000 ;
        RECT 505.120000 137.460000 506.320000 137.940000 ;
        RECT 505.120000 132.020000 506.320000 132.500000 ;
        RECT 545.600000 126.580000 546.800000 127.060000 ;
        RECT 545.600000 121.140000 546.800000 121.620000 ;
        RECT 545.600000 115.700000 546.800000 116.180000 ;
        RECT 545.600000 148.340000 546.800000 148.820000 ;
        RECT 545.600000 142.900000 546.800000 143.380000 ;
        RECT 545.600000 137.460000 546.800000 137.940000 ;
        RECT 545.600000 132.020000 546.800000 132.500000 ;
        RECT 415.120000 224.500000 416.320000 224.980000 ;
        RECT 370.120000 224.500000 371.320000 224.980000 ;
        RECT 325.120000 224.500000 326.320000 224.980000 ;
        RECT 280.120000 224.500000 281.320000 224.980000 ;
        RECT 280.120000 153.780000 281.320000 154.260000 ;
        RECT 280.120000 159.220000 281.320000 159.700000 ;
        RECT 280.120000 164.660000 281.320000 165.140000 ;
        RECT 280.120000 186.420000 281.320000 186.900000 ;
        RECT 280.120000 180.980000 281.320000 181.460000 ;
        RECT 280.120000 175.540000 281.320000 176.020000 ;
        RECT 280.120000 170.100000 281.320000 170.580000 ;
        RECT 325.120000 153.780000 326.320000 154.260000 ;
        RECT 325.120000 159.220000 326.320000 159.700000 ;
        RECT 325.120000 164.660000 326.320000 165.140000 ;
        RECT 325.120000 186.420000 326.320000 186.900000 ;
        RECT 325.120000 180.980000 326.320000 181.460000 ;
        RECT 325.120000 175.540000 326.320000 176.020000 ;
        RECT 325.120000 170.100000 326.320000 170.580000 ;
        RECT 280.120000 191.860000 281.320000 192.340000 ;
        RECT 280.120000 197.300000 281.320000 197.780000 ;
        RECT 280.120000 202.740000 281.320000 203.220000 ;
        RECT 280.120000 219.060000 281.320000 219.540000 ;
        RECT 280.120000 213.620000 281.320000 214.100000 ;
        RECT 280.120000 208.180000 281.320000 208.660000 ;
        RECT 325.120000 191.860000 326.320000 192.340000 ;
        RECT 325.120000 197.300000 326.320000 197.780000 ;
        RECT 325.120000 202.740000 326.320000 203.220000 ;
        RECT 325.120000 219.060000 326.320000 219.540000 ;
        RECT 325.120000 213.620000 326.320000 214.100000 ;
        RECT 325.120000 208.180000 326.320000 208.660000 ;
        RECT 370.120000 153.780000 371.320000 154.260000 ;
        RECT 370.120000 159.220000 371.320000 159.700000 ;
        RECT 370.120000 164.660000 371.320000 165.140000 ;
        RECT 370.120000 186.420000 371.320000 186.900000 ;
        RECT 370.120000 180.980000 371.320000 181.460000 ;
        RECT 370.120000 175.540000 371.320000 176.020000 ;
        RECT 370.120000 170.100000 371.320000 170.580000 ;
        RECT 415.120000 153.780000 416.320000 154.260000 ;
        RECT 415.120000 159.220000 416.320000 159.700000 ;
        RECT 415.120000 164.660000 416.320000 165.140000 ;
        RECT 415.120000 186.420000 416.320000 186.900000 ;
        RECT 415.120000 180.980000 416.320000 181.460000 ;
        RECT 415.120000 175.540000 416.320000 176.020000 ;
        RECT 415.120000 170.100000 416.320000 170.580000 ;
        RECT 370.120000 191.860000 371.320000 192.340000 ;
        RECT 370.120000 197.300000 371.320000 197.780000 ;
        RECT 370.120000 202.740000 371.320000 203.220000 ;
        RECT 370.120000 219.060000 371.320000 219.540000 ;
        RECT 370.120000 213.620000 371.320000 214.100000 ;
        RECT 370.120000 208.180000 371.320000 208.660000 ;
        RECT 415.120000 191.860000 416.320000 192.340000 ;
        RECT 415.120000 197.300000 416.320000 197.780000 ;
        RECT 415.120000 202.740000 416.320000 203.220000 ;
        RECT 415.120000 219.060000 416.320000 219.540000 ;
        RECT 415.120000 213.620000 416.320000 214.100000 ;
        RECT 415.120000 208.180000 416.320000 208.660000 ;
        RECT 280.120000 229.940000 281.320000 230.420000 ;
        RECT 280.120000 235.380000 281.320000 235.860000 ;
        RECT 280.120000 240.820000 281.320000 241.300000 ;
        RECT 280.120000 257.140000 281.320000 257.620000 ;
        RECT 280.120000 251.700000 281.320000 252.180000 ;
        RECT 280.120000 246.260000 281.320000 246.740000 ;
        RECT 325.120000 229.940000 326.320000 230.420000 ;
        RECT 325.120000 235.380000 326.320000 235.860000 ;
        RECT 325.120000 240.820000 326.320000 241.300000 ;
        RECT 325.120000 257.140000 326.320000 257.620000 ;
        RECT 325.120000 251.700000 326.320000 252.180000 ;
        RECT 325.120000 246.260000 326.320000 246.740000 ;
        RECT 280.120000 278.900000 281.320000 279.380000 ;
        RECT 280.120000 262.580000 281.320000 263.060000 ;
        RECT 280.120000 268.020000 281.320000 268.500000 ;
        RECT 280.120000 273.460000 281.320000 273.940000 ;
        RECT 280.120000 295.220000 281.320000 295.700000 ;
        RECT 280.120000 289.780000 281.320000 290.260000 ;
        RECT 280.120000 284.340000 281.320000 284.820000 ;
        RECT 325.120000 278.900000 326.320000 279.380000 ;
        RECT 325.120000 262.580000 326.320000 263.060000 ;
        RECT 325.120000 268.020000 326.320000 268.500000 ;
        RECT 325.120000 273.460000 326.320000 273.940000 ;
        RECT 325.120000 295.220000 326.320000 295.700000 ;
        RECT 325.120000 289.780000 326.320000 290.260000 ;
        RECT 325.120000 284.340000 326.320000 284.820000 ;
        RECT 370.120000 229.940000 371.320000 230.420000 ;
        RECT 370.120000 235.380000 371.320000 235.860000 ;
        RECT 370.120000 240.820000 371.320000 241.300000 ;
        RECT 370.120000 257.140000 371.320000 257.620000 ;
        RECT 370.120000 251.700000 371.320000 252.180000 ;
        RECT 370.120000 246.260000 371.320000 246.740000 ;
        RECT 415.120000 229.940000 416.320000 230.420000 ;
        RECT 415.120000 235.380000 416.320000 235.860000 ;
        RECT 415.120000 240.820000 416.320000 241.300000 ;
        RECT 415.120000 257.140000 416.320000 257.620000 ;
        RECT 415.120000 251.700000 416.320000 252.180000 ;
        RECT 415.120000 246.260000 416.320000 246.740000 ;
        RECT 370.120000 278.900000 371.320000 279.380000 ;
        RECT 370.120000 262.580000 371.320000 263.060000 ;
        RECT 370.120000 268.020000 371.320000 268.500000 ;
        RECT 370.120000 273.460000 371.320000 273.940000 ;
        RECT 370.120000 295.220000 371.320000 295.700000 ;
        RECT 370.120000 289.780000 371.320000 290.260000 ;
        RECT 370.120000 284.340000 371.320000 284.820000 ;
        RECT 415.120000 278.900000 416.320000 279.380000 ;
        RECT 415.120000 262.580000 416.320000 263.060000 ;
        RECT 415.120000 268.020000 416.320000 268.500000 ;
        RECT 415.120000 273.460000 416.320000 273.940000 ;
        RECT 415.120000 295.220000 416.320000 295.700000 ;
        RECT 415.120000 289.780000 416.320000 290.260000 ;
        RECT 415.120000 284.340000 416.320000 284.820000 ;
        RECT 545.600000 224.500000 546.800000 224.980000 ;
        RECT 505.120000 224.500000 506.320000 224.980000 ;
        RECT 460.120000 224.500000 461.320000 224.980000 ;
        RECT 460.120000 186.420000 461.320000 186.900000 ;
        RECT 460.120000 180.980000 461.320000 181.460000 ;
        RECT 460.120000 175.540000 461.320000 176.020000 ;
        RECT 460.120000 170.100000 461.320000 170.580000 ;
        RECT 460.120000 153.780000 461.320000 154.260000 ;
        RECT 460.120000 159.220000 461.320000 159.700000 ;
        RECT 460.120000 164.660000 461.320000 165.140000 ;
        RECT 460.120000 219.060000 461.320000 219.540000 ;
        RECT 460.120000 213.620000 461.320000 214.100000 ;
        RECT 460.120000 208.180000 461.320000 208.660000 ;
        RECT 460.120000 191.860000 461.320000 192.340000 ;
        RECT 460.120000 197.300000 461.320000 197.780000 ;
        RECT 460.120000 202.740000 461.320000 203.220000 ;
        RECT 505.120000 164.660000 506.320000 165.140000 ;
        RECT 505.120000 159.220000 506.320000 159.700000 ;
        RECT 505.120000 153.780000 506.320000 154.260000 ;
        RECT 505.120000 186.420000 506.320000 186.900000 ;
        RECT 505.120000 180.980000 506.320000 181.460000 ;
        RECT 505.120000 175.540000 506.320000 176.020000 ;
        RECT 505.120000 170.100000 506.320000 170.580000 ;
        RECT 545.600000 164.660000 546.800000 165.140000 ;
        RECT 545.600000 159.220000 546.800000 159.700000 ;
        RECT 545.600000 153.780000 546.800000 154.260000 ;
        RECT 545.600000 186.420000 546.800000 186.900000 ;
        RECT 545.600000 180.980000 546.800000 181.460000 ;
        RECT 545.600000 175.540000 546.800000 176.020000 ;
        RECT 545.600000 170.100000 546.800000 170.580000 ;
        RECT 505.120000 202.740000 506.320000 203.220000 ;
        RECT 505.120000 197.300000 506.320000 197.780000 ;
        RECT 505.120000 191.860000 506.320000 192.340000 ;
        RECT 505.120000 219.060000 506.320000 219.540000 ;
        RECT 505.120000 213.620000 506.320000 214.100000 ;
        RECT 505.120000 208.180000 506.320000 208.660000 ;
        RECT 545.600000 202.740000 546.800000 203.220000 ;
        RECT 545.600000 197.300000 546.800000 197.780000 ;
        RECT 545.600000 191.860000 546.800000 192.340000 ;
        RECT 545.600000 219.060000 546.800000 219.540000 ;
        RECT 545.600000 213.620000 546.800000 214.100000 ;
        RECT 545.600000 208.180000 546.800000 208.660000 ;
        RECT 460.120000 257.140000 461.320000 257.620000 ;
        RECT 460.120000 251.700000 461.320000 252.180000 ;
        RECT 460.120000 246.260000 461.320000 246.740000 ;
        RECT 460.120000 229.940000 461.320000 230.420000 ;
        RECT 460.120000 235.380000 461.320000 235.860000 ;
        RECT 460.120000 240.820000 461.320000 241.300000 ;
        RECT 460.120000 295.220000 461.320000 295.700000 ;
        RECT 460.120000 289.780000 461.320000 290.260000 ;
        RECT 460.120000 284.340000 461.320000 284.820000 ;
        RECT 460.120000 278.900000 461.320000 279.380000 ;
        RECT 460.120000 262.580000 461.320000 263.060000 ;
        RECT 460.120000 268.020000 461.320000 268.500000 ;
        RECT 460.120000 273.460000 461.320000 273.940000 ;
        RECT 505.120000 240.820000 506.320000 241.300000 ;
        RECT 505.120000 235.380000 506.320000 235.860000 ;
        RECT 505.120000 229.940000 506.320000 230.420000 ;
        RECT 505.120000 257.140000 506.320000 257.620000 ;
        RECT 505.120000 251.700000 506.320000 252.180000 ;
        RECT 505.120000 246.260000 506.320000 246.740000 ;
        RECT 545.600000 240.820000 546.800000 241.300000 ;
        RECT 545.600000 235.380000 546.800000 235.860000 ;
        RECT 545.600000 229.940000 546.800000 230.420000 ;
        RECT 545.600000 257.140000 546.800000 257.620000 ;
        RECT 545.600000 251.700000 546.800000 252.180000 ;
        RECT 545.600000 246.260000 546.800000 246.740000 ;
        RECT 505.120000 273.460000 506.320000 273.940000 ;
        RECT 505.120000 268.020000 506.320000 268.500000 ;
        RECT 505.120000 262.580000 506.320000 263.060000 ;
        RECT 505.120000 278.900000 506.320000 279.380000 ;
        RECT 505.120000 295.220000 506.320000 295.700000 ;
        RECT 505.120000 289.780000 506.320000 290.260000 ;
        RECT 505.120000 284.340000 506.320000 284.820000 ;
        RECT 545.600000 278.900000 546.800000 279.380000 ;
        RECT 545.600000 273.460000 546.800000 273.940000 ;
        RECT 545.600000 268.020000 546.800000 268.500000 ;
        RECT 545.600000 262.580000 546.800000 263.060000 ;
        RECT 545.600000 295.220000 546.800000 295.700000 ;
        RECT 545.600000 289.780000 546.800000 290.260000 ;
        RECT 545.600000 284.340000 546.800000 284.820000 ;
        RECT 3.360000 306.100000 4.560000 306.580000 ;
        RECT 9.955000 306.100000 11.320000 306.580000 ;
        RECT 3.360000 300.660000 4.560000 301.140000 ;
        RECT 9.955000 300.660000 11.320000 301.140000 ;
        RECT 3.360000 316.980000 4.560000 317.460000 ;
        RECT 9.955000 316.980000 11.320000 317.460000 ;
        RECT 3.360000 311.540000 4.560000 312.020000 ;
        RECT 9.955000 311.540000 11.320000 312.020000 ;
        RECT 3.360000 327.860000 4.560000 328.340000 ;
        RECT 9.955000 327.860000 11.320000 328.340000 ;
        RECT 3.360000 322.420000 4.560000 322.900000 ;
        RECT 9.955000 322.420000 11.320000 322.900000 ;
        RECT 3.360000 333.300000 4.560000 333.780000 ;
        RECT 9.955000 333.300000 11.320000 333.780000 ;
        RECT 3.360000 344.180000 4.560000 344.660000 ;
        RECT 9.955000 344.180000 11.320000 344.660000 ;
        RECT 3.360000 338.740000 4.560000 339.220000 ;
        RECT 9.955000 338.740000 11.320000 339.220000 ;
        RECT 3.360000 355.060000 4.560000 355.540000 ;
        RECT 9.955000 355.060000 11.320000 355.540000 ;
        RECT 3.360000 349.620000 4.560000 350.100000 ;
        RECT 9.955000 349.620000 11.320000 350.100000 ;
        RECT 3.360000 360.500000 4.560000 360.980000 ;
        RECT 9.955000 360.500000 11.320000 360.980000 ;
        RECT 3.360000 371.380000 4.560000 371.860000 ;
        RECT 9.955000 371.380000 11.320000 371.860000 ;
        RECT 3.360000 365.940000 4.560000 366.420000 ;
        RECT 9.955000 365.940000 11.320000 366.420000 ;
        RECT 55.120000 316.980000 56.320000 317.460000 ;
        RECT 55.120000 300.660000 56.320000 301.140000 ;
        RECT 55.120000 306.100000 56.320000 306.580000 ;
        RECT 55.120000 311.540000 56.320000 312.020000 ;
        RECT 55.120000 333.300000 56.320000 333.780000 ;
        RECT 55.120000 327.860000 56.320000 328.340000 ;
        RECT 55.120000 322.420000 56.320000 322.900000 ;
        RECT 100.120000 316.980000 101.320000 317.460000 ;
        RECT 100.120000 300.660000 101.320000 301.140000 ;
        RECT 100.120000 306.100000 101.320000 306.580000 ;
        RECT 100.120000 311.540000 101.320000 312.020000 ;
        RECT 100.120000 333.300000 101.320000 333.780000 ;
        RECT 100.120000 327.860000 101.320000 328.340000 ;
        RECT 100.120000 322.420000 101.320000 322.900000 ;
        RECT 55.120000 355.060000 56.320000 355.540000 ;
        RECT 55.120000 338.740000 56.320000 339.220000 ;
        RECT 55.120000 344.180000 56.320000 344.660000 ;
        RECT 55.120000 349.620000 56.320000 350.100000 ;
        RECT 55.120000 371.380000 56.320000 371.860000 ;
        RECT 55.120000 365.940000 56.320000 366.420000 ;
        RECT 55.120000 360.500000 56.320000 360.980000 ;
        RECT 100.120000 355.060000 101.320000 355.540000 ;
        RECT 100.120000 338.740000 101.320000 339.220000 ;
        RECT 100.120000 344.180000 101.320000 344.660000 ;
        RECT 100.120000 349.620000 101.320000 350.100000 ;
        RECT 100.120000 371.380000 101.320000 371.860000 ;
        RECT 100.120000 365.940000 101.320000 366.420000 ;
        RECT 100.120000 360.500000 101.320000 360.980000 ;
        RECT 3.360000 393.140000 4.560000 393.620000 ;
        RECT 9.955000 393.140000 11.320000 393.620000 ;
        RECT 3.360000 382.260000 4.560000 382.740000 ;
        RECT 9.955000 382.260000 11.320000 382.740000 ;
        RECT 3.360000 376.820000 4.560000 377.300000 ;
        RECT 9.955000 376.820000 11.320000 377.300000 ;
        RECT 3.360000 387.700000 4.560000 388.180000 ;
        RECT 9.955000 387.700000 11.320000 388.180000 ;
        RECT 3.360000 398.580000 4.560000 399.060000 ;
        RECT 9.955000 398.580000 11.320000 399.060000 ;
        RECT 3.360000 409.460000 4.560000 409.940000 ;
        RECT 3.360000 404.020000 4.560000 404.500000 ;
        RECT 9.955000 404.020000 11.320000 404.500000 ;
        RECT 9.955000 409.460000 11.320000 409.940000 ;
        RECT 3.360000 420.340000 4.560000 420.820000 ;
        RECT 9.955000 420.340000 11.320000 420.820000 ;
        RECT 3.360000 414.900000 4.560000 415.380000 ;
        RECT 9.955000 414.900000 11.320000 415.380000 ;
        RECT 3.360000 425.780000 4.560000 426.260000 ;
        RECT 9.955000 425.780000 11.320000 426.260000 ;
        RECT 3.360000 436.660000 4.560000 437.140000 ;
        RECT 9.955000 436.660000 11.320000 437.140000 ;
        RECT 3.360000 431.220000 4.560000 431.700000 ;
        RECT 9.955000 431.220000 11.320000 431.700000 ;
        RECT 3.360000 447.540000 4.560000 448.020000 ;
        RECT 9.955000 447.540000 11.320000 448.020000 ;
        RECT 3.360000 442.100000 4.560000 442.580000 ;
        RECT 9.955000 442.100000 11.320000 442.580000 ;
        RECT 55.120000 393.140000 56.320000 393.620000 ;
        RECT 55.120000 376.820000 56.320000 377.300000 ;
        RECT 55.120000 382.260000 56.320000 382.740000 ;
        RECT 55.120000 387.700000 56.320000 388.180000 ;
        RECT 55.120000 409.460000 56.320000 409.940000 ;
        RECT 55.120000 404.020000 56.320000 404.500000 ;
        RECT 55.120000 398.580000 56.320000 399.060000 ;
        RECT 100.120000 393.140000 101.320000 393.620000 ;
        RECT 100.120000 376.820000 101.320000 377.300000 ;
        RECT 100.120000 382.260000 101.320000 382.740000 ;
        RECT 100.120000 387.700000 101.320000 388.180000 ;
        RECT 100.120000 409.460000 101.320000 409.940000 ;
        RECT 100.120000 404.020000 101.320000 404.500000 ;
        RECT 100.120000 398.580000 101.320000 399.060000 ;
        RECT 55.120000 414.900000 56.320000 415.380000 ;
        RECT 55.120000 420.340000 56.320000 420.820000 ;
        RECT 55.120000 425.780000 56.320000 426.260000 ;
        RECT 55.120000 447.540000 56.320000 448.020000 ;
        RECT 55.120000 442.100000 56.320000 442.580000 ;
        RECT 55.120000 436.660000 56.320000 437.140000 ;
        RECT 55.120000 431.220000 56.320000 431.700000 ;
        RECT 100.120000 414.900000 101.320000 415.380000 ;
        RECT 100.120000 420.340000 101.320000 420.820000 ;
        RECT 100.120000 425.780000 101.320000 426.260000 ;
        RECT 100.120000 447.540000 101.320000 448.020000 ;
        RECT 100.120000 442.100000 101.320000 442.580000 ;
        RECT 100.120000 436.660000 101.320000 437.140000 ;
        RECT 100.120000 431.220000 101.320000 431.700000 ;
        RECT 145.120000 316.980000 146.320000 317.460000 ;
        RECT 145.120000 300.660000 146.320000 301.140000 ;
        RECT 145.120000 306.100000 146.320000 306.580000 ;
        RECT 145.120000 311.540000 146.320000 312.020000 ;
        RECT 145.120000 333.300000 146.320000 333.780000 ;
        RECT 145.120000 327.860000 146.320000 328.340000 ;
        RECT 145.120000 322.420000 146.320000 322.900000 ;
        RECT 190.120000 316.980000 191.320000 317.460000 ;
        RECT 190.120000 300.660000 191.320000 301.140000 ;
        RECT 190.120000 306.100000 191.320000 306.580000 ;
        RECT 190.120000 311.540000 191.320000 312.020000 ;
        RECT 190.120000 333.300000 191.320000 333.780000 ;
        RECT 190.120000 327.860000 191.320000 328.340000 ;
        RECT 190.120000 322.420000 191.320000 322.900000 ;
        RECT 145.120000 355.060000 146.320000 355.540000 ;
        RECT 145.120000 338.740000 146.320000 339.220000 ;
        RECT 145.120000 344.180000 146.320000 344.660000 ;
        RECT 145.120000 349.620000 146.320000 350.100000 ;
        RECT 145.120000 371.380000 146.320000 371.860000 ;
        RECT 145.120000 365.940000 146.320000 366.420000 ;
        RECT 145.120000 360.500000 146.320000 360.980000 ;
        RECT 190.120000 355.060000 191.320000 355.540000 ;
        RECT 190.120000 338.740000 191.320000 339.220000 ;
        RECT 190.120000 344.180000 191.320000 344.660000 ;
        RECT 190.120000 349.620000 191.320000 350.100000 ;
        RECT 190.120000 371.380000 191.320000 371.860000 ;
        RECT 190.120000 365.940000 191.320000 366.420000 ;
        RECT 190.120000 360.500000 191.320000 360.980000 ;
        RECT 235.120000 333.300000 236.320000 333.780000 ;
        RECT 235.120000 327.860000 236.320000 328.340000 ;
        RECT 235.120000 322.420000 236.320000 322.900000 ;
        RECT 235.120000 316.980000 236.320000 317.460000 ;
        RECT 235.120000 300.660000 236.320000 301.140000 ;
        RECT 235.120000 306.100000 236.320000 306.580000 ;
        RECT 235.120000 311.540000 236.320000 312.020000 ;
        RECT 235.120000 371.380000 236.320000 371.860000 ;
        RECT 235.120000 365.940000 236.320000 366.420000 ;
        RECT 235.120000 360.500000 236.320000 360.980000 ;
        RECT 235.120000 355.060000 236.320000 355.540000 ;
        RECT 235.120000 338.740000 236.320000 339.220000 ;
        RECT 235.120000 344.180000 236.320000 344.660000 ;
        RECT 235.120000 349.620000 236.320000 350.100000 ;
        RECT 145.120000 393.140000 146.320000 393.620000 ;
        RECT 145.120000 376.820000 146.320000 377.300000 ;
        RECT 145.120000 382.260000 146.320000 382.740000 ;
        RECT 145.120000 387.700000 146.320000 388.180000 ;
        RECT 145.120000 409.460000 146.320000 409.940000 ;
        RECT 145.120000 404.020000 146.320000 404.500000 ;
        RECT 145.120000 398.580000 146.320000 399.060000 ;
        RECT 190.120000 393.140000 191.320000 393.620000 ;
        RECT 190.120000 376.820000 191.320000 377.300000 ;
        RECT 190.120000 382.260000 191.320000 382.740000 ;
        RECT 190.120000 387.700000 191.320000 388.180000 ;
        RECT 190.120000 409.460000 191.320000 409.940000 ;
        RECT 190.120000 404.020000 191.320000 404.500000 ;
        RECT 190.120000 398.580000 191.320000 399.060000 ;
        RECT 145.120000 414.900000 146.320000 415.380000 ;
        RECT 145.120000 420.340000 146.320000 420.820000 ;
        RECT 145.120000 425.780000 146.320000 426.260000 ;
        RECT 145.120000 447.540000 146.320000 448.020000 ;
        RECT 145.120000 442.100000 146.320000 442.580000 ;
        RECT 145.120000 436.660000 146.320000 437.140000 ;
        RECT 145.120000 431.220000 146.320000 431.700000 ;
        RECT 190.120000 414.900000 191.320000 415.380000 ;
        RECT 190.120000 420.340000 191.320000 420.820000 ;
        RECT 190.120000 425.780000 191.320000 426.260000 ;
        RECT 190.120000 447.540000 191.320000 448.020000 ;
        RECT 190.120000 442.100000 191.320000 442.580000 ;
        RECT 190.120000 436.660000 191.320000 437.140000 ;
        RECT 190.120000 431.220000 191.320000 431.700000 ;
        RECT 235.120000 409.460000 236.320000 409.940000 ;
        RECT 235.120000 404.020000 236.320000 404.500000 ;
        RECT 235.120000 398.580000 236.320000 399.060000 ;
        RECT 235.120000 376.820000 236.320000 377.300000 ;
        RECT 235.120000 382.260000 236.320000 382.740000 ;
        RECT 235.120000 387.700000 236.320000 388.180000 ;
        RECT 235.120000 393.140000 236.320000 393.620000 ;
        RECT 235.120000 447.540000 236.320000 448.020000 ;
        RECT 235.120000 442.100000 236.320000 442.580000 ;
        RECT 235.120000 436.660000 236.320000 437.140000 ;
        RECT 235.120000 414.900000 236.320000 415.380000 ;
        RECT 235.120000 420.340000 236.320000 420.820000 ;
        RECT 235.120000 425.780000 236.320000 426.260000 ;
        RECT 235.120000 431.220000 236.320000 431.700000 ;
        RECT 3.360000 458.420000 4.560000 458.900000 ;
        RECT 3.360000 452.980000 4.560000 453.460000 ;
        RECT 9.955000 452.980000 11.320000 453.460000 ;
        RECT 9.955000 458.420000 11.320000 458.900000 ;
        RECT 3.360000 463.860000 4.560000 464.340000 ;
        RECT 9.955000 463.860000 11.320000 464.340000 ;
        RECT 3.360000 474.740000 4.560000 475.220000 ;
        RECT 9.955000 474.740000 11.320000 475.220000 ;
        RECT 3.360000 469.300000 4.560000 469.780000 ;
        RECT 9.955000 469.300000 11.320000 469.780000 ;
        RECT 3.360000 485.620000 4.560000 486.100000 ;
        RECT 9.955000 485.620000 11.320000 486.100000 ;
        RECT 3.360000 480.180000 4.560000 480.660000 ;
        RECT 9.955000 480.180000 11.320000 480.660000 ;
        RECT 3.360000 496.500000 4.560000 496.980000 ;
        RECT 9.955000 496.500000 11.320000 496.980000 ;
        RECT 3.360000 491.060000 4.560000 491.540000 ;
        RECT 9.955000 491.060000 11.320000 491.540000 ;
        RECT 3.360000 501.940000 4.560000 502.420000 ;
        RECT 9.955000 501.940000 11.320000 502.420000 ;
        RECT 3.360000 512.820000 4.560000 513.300000 ;
        RECT 9.955000 512.820000 11.320000 513.300000 ;
        RECT 3.360000 507.380000 4.560000 507.860000 ;
        RECT 9.955000 507.380000 11.320000 507.860000 ;
        RECT 3.360000 523.700000 4.560000 524.180000 ;
        RECT 9.955000 523.700000 11.320000 524.180000 ;
        RECT 3.360000 518.260000 4.560000 518.740000 ;
        RECT 9.955000 518.260000 11.320000 518.740000 ;
        RECT 55.120000 452.980000 56.320000 453.460000 ;
        RECT 55.120000 458.420000 56.320000 458.900000 ;
        RECT 55.120000 463.860000 56.320000 464.340000 ;
        RECT 55.120000 485.620000 56.320000 486.100000 ;
        RECT 55.120000 480.180000 56.320000 480.660000 ;
        RECT 55.120000 474.740000 56.320000 475.220000 ;
        RECT 55.120000 469.300000 56.320000 469.780000 ;
        RECT 100.120000 452.980000 101.320000 453.460000 ;
        RECT 100.120000 458.420000 101.320000 458.900000 ;
        RECT 100.120000 463.860000 101.320000 464.340000 ;
        RECT 100.120000 485.620000 101.320000 486.100000 ;
        RECT 100.120000 480.180000 101.320000 480.660000 ;
        RECT 100.120000 474.740000 101.320000 475.220000 ;
        RECT 100.120000 469.300000 101.320000 469.780000 ;
        RECT 55.120000 491.060000 56.320000 491.540000 ;
        RECT 55.120000 496.500000 56.320000 496.980000 ;
        RECT 55.120000 501.940000 56.320000 502.420000 ;
        RECT 55.120000 523.700000 56.320000 524.180000 ;
        RECT 55.120000 518.260000 56.320000 518.740000 ;
        RECT 55.120000 512.820000 56.320000 513.300000 ;
        RECT 55.120000 507.380000 56.320000 507.860000 ;
        RECT 100.120000 491.060000 101.320000 491.540000 ;
        RECT 100.120000 496.500000 101.320000 496.980000 ;
        RECT 100.120000 501.940000 101.320000 502.420000 ;
        RECT 100.120000 523.700000 101.320000 524.180000 ;
        RECT 100.120000 518.260000 101.320000 518.740000 ;
        RECT 100.120000 512.820000 101.320000 513.300000 ;
        RECT 100.120000 507.380000 101.320000 507.860000 ;
        RECT 3.360000 529.140000 4.560000 529.620000 ;
        RECT 9.955000 529.140000 11.320000 529.620000 ;
        RECT 3.360000 540.020000 4.560000 540.500000 ;
        RECT 9.955000 540.020000 11.320000 540.500000 ;
        RECT 3.360000 534.580000 4.560000 535.060000 ;
        RECT 9.955000 534.580000 11.320000 535.060000 ;
        RECT 3.360000 550.900000 4.560000 551.380000 ;
        RECT 9.955000 550.900000 11.320000 551.380000 ;
        RECT 3.360000 545.460000 4.560000 545.940000 ;
        RECT 9.955000 545.460000 11.320000 545.940000 ;
        RECT 3.360000 561.780000 4.560000 562.260000 ;
        RECT 9.955000 561.780000 11.320000 562.260000 ;
        RECT 3.360000 556.340000 4.560000 556.820000 ;
        RECT 9.955000 556.340000 11.320000 556.820000 ;
        RECT 3.360000 567.220000 4.560000 567.700000 ;
        RECT 9.955000 567.220000 11.320000 567.700000 ;
        RECT 3.360000 578.100000 4.560000 578.580000 ;
        RECT 3.360000 572.660000 4.560000 573.140000 ;
        RECT 9.955000 572.660000 11.320000 573.140000 ;
        RECT 9.955000 578.100000 11.320000 578.580000 ;
        RECT 3.360000 588.980000 4.560000 589.460000 ;
        RECT 9.955000 588.980000 11.320000 589.460000 ;
        RECT 3.360000 583.540000 4.560000 584.020000 ;
        RECT 9.955000 583.540000 11.320000 584.020000 ;
        RECT 55.120000 529.140000 56.320000 529.620000 ;
        RECT 55.120000 534.580000 56.320000 535.060000 ;
        RECT 55.120000 540.020000 56.320000 540.500000 ;
        RECT 55.120000 561.780000 56.320000 562.260000 ;
        RECT 55.120000 556.340000 56.320000 556.820000 ;
        RECT 55.120000 550.900000 56.320000 551.380000 ;
        RECT 55.120000 545.460000 56.320000 545.940000 ;
        RECT 100.120000 529.140000 101.320000 529.620000 ;
        RECT 100.120000 534.580000 101.320000 535.060000 ;
        RECT 100.120000 540.020000 101.320000 540.500000 ;
        RECT 100.120000 561.780000 101.320000 562.260000 ;
        RECT 100.120000 556.340000 101.320000 556.820000 ;
        RECT 100.120000 550.900000 101.320000 551.380000 ;
        RECT 100.120000 545.460000 101.320000 545.940000 ;
        RECT 55.120000 567.220000 56.320000 567.700000 ;
        RECT 55.120000 572.660000 56.320000 573.140000 ;
        RECT 55.120000 578.100000 56.320000 578.580000 ;
        RECT 55.120000 583.540000 56.320000 584.020000 ;
        RECT 55.120000 588.980000 56.320000 589.460000 ;
        RECT 100.120000 567.220000 101.320000 567.700000 ;
        RECT 100.120000 572.660000 101.320000 573.140000 ;
        RECT 100.120000 578.100000 101.320000 578.580000 ;
        RECT 100.120000 583.540000 101.320000 584.020000 ;
        RECT 100.120000 588.980000 101.320000 589.460000 ;
        RECT 145.120000 452.980000 146.320000 453.460000 ;
        RECT 145.120000 458.420000 146.320000 458.900000 ;
        RECT 145.120000 463.860000 146.320000 464.340000 ;
        RECT 145.120000 485.620000 146.320000 486.100000 ;
        RECT 145.120000 480.180000 146.320000 480.660000 ;
        RECT 145.120000 474.740000 146.320000 475.220000 ;
        RECT 145.120000 469.300000 146.320000 469.780000 ;
        RECT 190.120000 452.980000 191.320000 453.460000 ;
        RECT 190.120000 458.420000 191.320000 458.900000 ;
        RECT 190.120000 463.860000 191.320000 464.340000 ;
        RECT 190.120000 485.620000 191.320000 486.100000 ;
        RECT 190.120000 480.180000 191.320000 480.660000 ;
        RECT 190.120000 474.740000 191.320000 475.220000 ;
        RECT 190.120000 469.300000 191.320000 469.780000 ;
        RECT 145.120000 491.060000 146.320000 491.540000 ;
        RECT 145.120000 496.500000 146.320000 496.980000 ;
        RECT 145.120000 501.940000 146.320000 502.420000 ;
        RECT 145.120000 523.700000 146.320000 524.180000 ;
        RECT 145.120000 518.260000 146.320000 518.740000 ;
        RECT 145.120000 512.820000 146.320000 513.300000 ;
        RECT 145.120000 507.380000 146.320000 507.860000 ;
        RECT 190.120000 491.060000 191.320000 491.540000 ;
        RECT 190.120000 496.500000 191.320000 496.980000 ;
        RECT 190.120000 501.940000 191.320000 502.420000 ;
        RECT 190.120000 523.700000 191.320000 524.180000 ;
        RECT 190.120000 518.260000 191.320000 518.740000 ;
        RECT 190.120000 512.820000 191.320000 513.300000 ;
        RECT 190.120000 507.380000 191.320000 507.860000 ;
        RECT 235.120000 485.620000 236.320000 486.100000 ;
        RECT 235.120000 480.180000 236.320000 480.660000 ;
        RECT 235.120000 474.740000 236.320000 475.220000 ;
        RECT 235.120000 469.300000 236.320000 469.780000 ;
        RECT 235.120000 452.980000 236.320000 453.460000 ;
        RECT 235.120000 458.420000 236.320000 458.900000 ;
        RECT 235.120000 463.860000 236.320000 464.340000 ;
        RECT 235.120000 523.700000 236.320000 524.180000 ;
        RECT 235.120000 518.260000 236.320000 518.740000 ;
        RECT 235.120000 512.820000 236.320000 513.300000 ;
        RECT 235.120000 507.380000 236.320000 507.860000 ;
        RECT 235.120000 491.060000 236.320000 491.540000 ;
        RECT 235.120000 496.500000 236.320000 496.980000 ;
        RECT 235.120000 501.940000 236.320000 502.420000 ;
        RECT 145.120000 529.140000 146.320000 529.620000 ;
        RECT 145.120000 534.580000 146.320000 535.060000 ;
        RECT 145.120000 540.020000 146.320000 540.500000 ;
        RECT 145.120000 561.780000 146.320000 562.260000 ;
        RECT 145.120000 556.340000 146.320000 556.820000 ;
        RECT 145.120000 550.900000 146.320000 551.380000 ;
        RECT 145.120000 545.460000 146.320000 545.940000 ;
        RECT 190.120000 529.140000 191.320000 529.620000 ;
        RECT 190.120000 534.580000 191.320000 535.060000 ;
        RECT 190.120000 540.020000 191.320000 540.500000 ;
        RECT 190.120000 561.780000 191.320000 562.260000 ;
        RECT 190.120000 556.340000 191.320000 556.820000 ;
        RECT 190.120000 550.900000 191.320000 551.380000 ;
        RECT 190.120000 545.460000 191.320000 545.940000 ;
        RECT 145.120000 567.220000 146.320000 567.700000 ;
        RECT 145.120000 572.660000 146.320000 573.140000 ;
        RECT 145.120000 578.100000 146.320000 578.580000 ;
        RECT 145.120000 583.540000 146.320000 584.020000 ;
        RECT 145.120000 588.980000 146.320000 589.460000 ;
        RECT 190.120000 567.220000 191.320000 567.700000 ;
        RECT 190.120000 572.660000 191.320000 573.140000 ;
        RECT 190.120000 578.100000 191.320000 578.580000 ;
        RECT 190.120000 583.540000 191.320000 584.020000 ;
        RECT 190.120000 588.980000 191.320000 589.460000 ;
        RECT 235.120000 561.780000 236.320000 562.260000 ;
        RECT 235.120000 556.340000 236.320000 556.820000 ;
        RECT 235.120000 550.900000 236.320000 551.380000 ;
        RECT 235.120000 545.460000 236.320000 545.940000 ;
        RECT 235.120000 529.140000 236.320000 529.620000 ;
        RECT 235.120000 534.580000 236.320000 535.060000 ;
        RECT 235.120000 540.020000 236.320000 540.500000 ;
        RECT 235.120000 567.220000 236.320000 567.700000 ;
        RECT 235.120000 572.660000 236.320000 573.140000 ;
        RECT 235.120000 578.100000 236.320000 578.580000 ;
        RECT 235.120000 583.540000 236.320000 584.020000 ;
        RECT 235.120000 588.980000 236.320000 589.460000 ;
        RECT 280.120000 316.980000 281.320000 317.460000 ;
        RECT 280.120000 300.660000 281.320000 301.140000 ;
        RECT 280.120000 306.100000 281.320000 306.580000 ;
        RECT 280.120000 311.540000 281.320000 312.020000 ;
        RECT 280.120000 333.300000 281.320000 333.780000 ;
        RECT 280.120000 327.860000 281.320000 328.340000 ;
        RECT 280.120000 322.420000 281.320000 322.900000 ;
        RECT 325.120000 316.980000 326.320000 317.460000 ;
        RECT 325.120000 300.660000 326.320000 301.140000 ;
        RECT 325.120000 306.100000 326.320000 306.580000 ;
        RECT 325.120000 311.540000 326.320000 312.020000 ;
        RECT 325.120000 333.300000 326.320000 333.780000 ;
        RECT 325.120000 327.860000 326.320000 328.340000 ;
        RECT 325.120000 322.420000 326.320000 322.900000 ;
        RECT 280.120000 355.060000 281.320000 355.540000 ;
        RECT 280.120000 338.740000 281.320000 339.220000 ;
        RECT 280.120000 344.180000 281.320000 344.660000 ;
        RECT 280.120000 349.620000 281.320000 350.100000 ;
        RECT 280.120000 371.380000 281.320000 371.860000 ;
        RECT 280.120000 365.940000 281.320000 366.420000 ;
        RECT 280.120000 360.500000 281.320000 360.980000 ;
        RECT 325.120000 355.060000 326.320000 355.540000 ;
        RECT 325.120000 338.740000 326.320000 339.220000 ;
        RECT 325.120000 344.180000 326.320000 344.660000 ;
        RECT 325.120000 349.620000 326.320000 350.100000 ;
        RECT 325.120000 371.380000 326.320000 371.860000 ;
        RECT 325.120000 365.940000 326.320000 366.420000 ;
        RECT 325.120000 360.500000 326.320000 360.980000 ;
        RECT 370.120000 316.980000 371.320000 317.460000 ;
        RECT 370.120000 300.660000 371.320000 301.140000 ;
        RECT 370.120000 306.100000 371.320000 306.580000 ;
        RECT 370.120000 311.540000 371.320000 312.020000 ;
        RECT 370.120000 333.300000 371.320000 333.780000 ;
        RECT 370.120000 327.860000 371.320000 328.340000 ;
        RECT 370.120000 322.420000 371.320000 322.900000 ;
        RECT 415.120000 316.980000 416.320000 317.460000 ;
        RECT 415.120000 300.660000 416.320000 301.140000 ;
        RECT 415.120000 306.100000 416.320000 306.580000 ;
        RECT 415.120000 311.540000 416.320000 312.020000 ;
        RECT 415.120000 333.300000 416.320000 333.780000 ;
        RECT 415.120000 327.860000 416.320000 328.340000 ;
        RECT 415.120000 322.420000 416.320000 322.900000 ;
        RECT 370.120000 355.060000 371.320000 355.540000 ;
        RECT 370.120000 338.740000 371.320000 339.220000 ;
        RECT 370.120000 344.180000 371.320000 344.660000 ;
        RECT 370.120000 349.620000 371.320000 350.100000 ;
        RECT 370.120000 371.380000 371.320000 371.860000 ;
        RECT 370.120000 365.940000 371.320000 366.420000 ;
        RECT 370.120000 360.500000 371.320000 360.980000 ;
        RECT 415.120000 355.060000 416.320000 355.540000 ;
        RECT 415.120000 338.740000 416.320000 339.220000 ;
        RECT 415.120000 344.180000 416.320000 344.660000 ;
        RECT 415.120000 349.620000 416.320000 350.100000 ;
        RECT 415.120000 371.380000 416.320000 371.860000 ;
        RECT 415.120000 365.940000 416.320000 366.420000 ;
        RECT 415.120000 360.500000 416.320000 360.980000 ;
        RECT 280.120000 393.140000 281.320000 393.620000 ;
        RECT 280.120000 376.820000 281.320000 377.300000 ;
        RECT 280.120000 382.260000 281.320000 382.740000 ;
        RECT 280.120000 387.700000 281.320000 388.180000 ;
        RECT 280.120000 409.460000 281.320000 409.940000 ;
        RECT 280.120000 404.020000 281.320000 404.500000 ;
        RECT 280.120000 398.580000 281.320000 399.060000 ;
        RECT 325.120000 393.140000 326.320000 393.620000 ;
        RECT 325.120000 376.820000 326.320000 377.300000 ;
        RECT 325.120000 382.260000 326.320000 382.740000 ;
        RECT 325.120000 387.700000 326.320000 388.180000 ;
        RECT 325.120000 409.460000 326.320000 409.940000 ;
        RECT 325.120000 404.020000 326.320000 404.500000 ;
        RECT 325.120000 398.580000 326.320000 399.060000 ;
        RECT 280.120000 414.900000 281.320000 415.380000 ;
        RECT 280.120000 420.340000 281.320000 420.820000 ;
        RECT 280.120000 425.780000 281.320000 426.260000 ;
        RECT 280.120000 447.540000 281.320000 448.020000 ;
        RECT 280.120000 442.100000 281.320000 442.580000 ;
        RECT 280.120000 436.660000 281.320000 437.140000 ;
        RECT 280.120000 431.220000 281.320000 431.700000 ;
        RECT 325.120000 414.900000 326.320000 415.380000 ;
        RECT 325.120000 420.340000 326.320000 420.820000 ;
        RECT 325.120000 425.780000 326.320000 426.260000 ;
        RECT 325.120000 447.540000 326.320000 448.020000 ;
        RECT 325.120000 442.100000 326.320000 442.580000 ;
        RECT 325.120000 436.660000 326.320000 437.140000 ;
        RECT 325.120000 431.220000 326.320000 431.700000 ;
        RECT 370.120000 393.140000 371.320000 393.620000 ;
        RECT 370.120000 376.820000 371.320000 377.300000 ;
        RECT 370.120000 382.260000 371.320000 382.740000 ;
        RECT 370.120000 387.700000 371.320000 388.180000 ;
        RECT 370.120000 409.460000 371.320000 409.940000 ;
        RECT 370.120000 404.020000 371.320000 404.500000 ;
        RECT 370.120000 398.580000 371.320000 399.060000 ;
        RECT 415.120000 393.140000 416.320000 393.620000 ;
        RECT 415.120000 376.820000 416.320000 377.300000 ;
        RECT 415.120000 382.260000 416.320000 382.740000 ;
        RECT 415.120000 387.700000 416.320000 388.180000 ;
        RECT 415.120000 409.460000 416.320000 409.940000 ;
        RECT 415.120000 404.020000 416.320000 404.500000 ;
        RECT 415.120000 398.580000 416.320000 399.060000 ;
        RECT 370.120000 414.900000 371.320000 415.380000 ;
        RECT 370.120000 420.340000 371.320000 420.820000 ;
        RECT 370.120000 425.780000 371.320000 426.260000 ;
        RECT 370.120000 447.540000 371.320000 448.020000 ;
        RECT 370.120000 442.100000 371.320000 442.580000 ;
        RECT 370.120000 436.660000 371.320000 437.140000 ;
        RECT 370.120000 431.220000 371.320000 431.700000 ;
        RECT 415.120000 414.900000 416.320000 415.380000 ;
        RECT 415.120000 420.340000 416.320000 420.820000 ;
        RECT 415.120000 425.780000 416.320000 426.260000 ;
        RECT 415.120000 447.540000 416.320000 448.020000 ;
        RECT 415.120000 442.100000 416.320000 442.580000 ;
        RECT 415.120000 436.660000 416.320000 437.140000 ;
        RECT 415.120000 431.220000 416.320000 431.700000 ;
        RECT 460.120000 333.300000 461.320000 333.780000 ;
        RECT 460.120000 327.860000 461.320000 328.340000 ;
        RECT 460.120000 322.420000 461.320000 322.900000 ;
        RECT 460.120000 316.980000 461.320000 317.460000 ;
        RECT 460.120000 300.660000 461.320000 301.140000 ;
        RECT 460.120000 306.100000 461.320000 306.580000 ;
        RECT 460.120000 311.540000 461.320000 312.020000 ;
        RECT 460.120000 371.380000 461.320000 371.860000 ;
        RECT 460.120000 365.940000 461.320000 366.420000 ;
        RECT 460.120000 360.500000 461.320000 360.980000 ;
        RECT 460.120000 355.060000 461.320000 355.540000 ;
        RECT 460.120000 338.740000 461.320000 339.220000 ;
        RECT 460.120000 344.180000 461.320000 344.660000 ;
        RECT 460.120000 349.620000 461.320000 350.100000 ;
        RECT 505.120000 311.540000 506.320000 312.020000 ;
        RECT 505.120000 306.100000 506.320000 306.580000 ;
        RECT 505.120000 300.660000 506.320000 301.140000 ;
        RECT 505.120000 316.980000 506.320000 317.460000 ;
        RECT 505.120000 333.300000 506.320000 333.780000 ;
        RECT 505.120000 327.860000 506.320000 328.340000 ;
        RECT 505.120000 322.420000 506.320000 322.900000 ;
        RECT 545.600000 316.980000 546.800000 317.460000 ;
        RECT 545.600000 311.540000 546.800000 312.020000 ;
        RECT 545.600000 306.100000 546.800000 306.580000 ;
        RECT 545.600000 300.660000 546.800000 301.140000 ;
        RECT 545.600000 333.300000 546.800000 333.780000 ;
        RECT 545.600000 327.860000 546.800000 328.340000 ;
        RECT 545.600000 322.420000 546.800000 322.900000 ;
        RECT 505.120000 349.620000 506.320000 350.100000 ;
        RECT 505.120000 344.180000 506.320000 344.660000 ;
        RECT 505.120000 338.740000 506.320000 339.220000 ;
        RECT 505.120000 355.060000 506.320000 355.540000 ;
        RECT 505.120000 371.380000 506.320000 371.860000 ;
        RECT 505.120000 365.940000 506.320000 366.420000 ;
        RECT 505.120000 360.500000 506.320000 360.980000 ;
        RECT 545.600000 355.060000 546.800000 355.540000 ;
        RECT 545.600000 349.620000 546.800000 350.100000 ;
        RECT 545.600000 344.180000 546.800000 344.660000 ;
        RECT 545.600000 338.740000 546.800000 339.220000 ;
        RECT 545.600000 371.380000 546.800000 371.860000 ;
        RECT 545.600000 365.940000 546.800000 366.420000 ;
        RECT 545.600000 360.500000 546.800000 360.980000 ;
        RECT 460.120000 409.460000 461.320000 409.940000 ;
        RECT 460.120000 404.020000 461.320000 404.500000 ;
        RECT 460.120000 398.580000 461.320000 399.060000 ;
        RECT 460.120000 376.820000 461.320000 377.300000 ;
        RECT 460.120000 382.260000 461.320000 382.740000 ;
        RECT 460.120000 387.700000 461.320000 388.180000 ;
        RECT 460.120000 393.140000 461.320000 393.620000 ;
        RECT 460.120000 447.540000 461.320000 448.020000 ;
        RECT 460.120000 442.100000 461.320000 442.580000 ;
        RECT 460.120000 436.660000 461.320000 437.140000 ;
        RECT 460.120000 414.900000 461.320000 415.380000 ;
        RECT 460.120000 420.340000 461.320000 420.820000 ;
        RECT 460.120000 425.780000 461.320000 426.260000 ;
        RECT 460.120000 431.220000 461.320000 431.700000 ;
        RECT 505.120000 393.140000 506.320000 393.620000 ;
        RECT 505.120000 387.700000 506.320000 388.180000 ;
        RECT 505.120000 382.260000 506.320000 382.740000 ;
        RECT 505.120000 376.820000 506.320000 377.300000 ;
        RECT 505.120000 409.460000 506.320000 409.940000 ;
        RECT 505.120000 404.020000 506.320000 404.500000 ;
        RECT 505.120000 398.580000 506.320000 399.060000 ;
        RECT 545.600000 393.140000 546.800000 393.620000 ;
        RECT 545.600000 387.700000 546.800000 388.180000 ;
        RECT 545.600000 376.820000 546.800000 377.300000 ;
        RECT 545.600000 382.260000 546.800000 382.740000 ;
        RECT 545.600000 409.460000 546.800000 409.940000 ;
        RECT 545.600000 404.020000 546.800000 404.500000 ;
        RECT 545.600000 398.580000 546.800000 399.060000 ;
        RECT 505.120000 425.780000 506.320000 426.260000 ;
        RECT 505.120000 420.340000 506.320000 420.820000 ;
        RECT 505.120000 414.900000 506.320000 415.380000 ;
        RECT 505.120000 447.540000 506.320000 448.020000 ;
        RECT 505.120000 442.100000 506.320000 442.580000 ;
        RECT 505.120000 431.220000 506.320000 431.700000 ;
        RECT 505.120000 436.660000 506.320000 437.140000 ;
        RECT 545.600000 425.780000 546.800000 426.260000 ;
        RECT 545.600000 414.900000 546.800000 415.380000 ;
        RECT 545.600000 420.340000 546.800000 420.820000 ;
        RECT 545.600000 447.540000 546.800000 448.020000 ;
        RECT 545.600000 442.100000 546.800000 442.580000 ;
        RECT 545.600000 436.660000 546.800000 437.140000 ;
        RECT 545.600000 431.220000 546.800000 431.700000 ;
        RECT 280.120000 452.980000 281.320000 453.460000 ;
        RECT 280.120000 458.420000 281.320000 458.900000 ;
        RECT 280.120000 463.860000 281.320000 464.340000 ;
        RECT 280.120000 485.620000 281.320000 486.100000 ;
        RECT 280.120000 480.180000 281.320000 480.660000 ;
        RECT 280.120000 474.740000 281.320000 475.220000 ;
        RECT 280.120000 469.300000 281.320000 469.780000 ;
        RECT 325.120000 452.980000 326.320000 453.460000 ;
        RECT 325.120000 458.420000 326.320000 458.900000 ;
        RECT 325.120000 463.860000 326.320000 464.340000 ;
        RECT 325.120000 485.620000 326.320000 486.100000 ;
        RECT 325.120000 480.180000 326.320000 480.660000 ;
        RECT 325.120000 474.740000 326.320000 475.220000 ;
        RECT 325.120000 469.300000 326.320000 469.780000 ;
        RECT 280.120000 491.060000 281.320000 491.540000 ;
        RECT 280.120000 496.500000 281.320000 496.980000 ;
        RECT 280.120000 501.940000 281.320000 502.420000 ;
        RECT 280.120000 523.700000 281.320000 524.180000 ;
        RECT 280.120000 518.260000 281.320000 518.740000 ;
        RECT 280.120000 512.820000 281.320000 513.300000 ;
        RECT 280.120000 507.380000 281.320000 507.860000 ;
        RECT 325.120000 491.060000 326.320000 491.540000 ;
        RECT 325.120000 496.500000 326.320000 496.980000 ;
        RECT 325.120000 501.940000 326.320000 502.420000 ;
        RECT 325.120000 523.700000 326.320000 524.180000 ;
        RECT 325.120000 518.260000 326.320000 518.740000 ;
        RECT 325.120000 512.820000 326.320000 513.300000 ;
        RECT 325.120000 507.380000 326.320000 507.860000 ;
        RECT 370.120000 452.980000 371.320000 453.460000 ;
        RECT 370.120000 458.420000 371.320000 458.900000 ;
        RECT 370.120000 463.860000 371.320000 464.340000 ;
        RECT 370.120000 485.620000 371.320000 486.100000 ;
        RECT 370.120000 480.180000 371.320000 480.660000 ;
        RECT 370.120000 474.740000 371.320000 475.220000 ;
        RECT 370.120000 469.300000 371.320000 469.780000 ;
        RECT 415.120000 452.980000 416.320000 453.460000 ;
        RECT 415.120000 458.420000 416.320000 458.900000 ;
        RECT 415.120000 463.860000 416.320000 464.340000 ;
        RECT 415.120000 485.620000 416.320000 486.100000 ;
        RECT 415.120000 480.180000 416.320000 480.660000 ;
        RECT 415.120000 474.740000 416.320000 475.220000 ;
        RECT 415.120000 469.300000 416.320000 469.780000 ;
        RECT 370.120000 491.060000 371.320000 491.540000 ;
        RECT 370.120000 496.500000 371.320000 496.980000 ;
        RECT 370.120000 501.940000 371.320000 502.420000 ;
        RECT 370.120000 523.700000 371.320000 524.180000 ;
        RECT 370.120000 518.260000 371.320000 518.740000 ;
        RECT 370.120000 512.820000 371.320000 513.300000 ;
        RECT 370.120000 507.380000 371.320000 507.860000 ;
        RECT 415.120000 491.060000 416.320000 491.540000 ;
        RECT 415.120000 496.500000 416.320000 496.980000 ;
        RECT 415.120000 501.940000 416.320000 502.420000 ;
        RECT 415.120000 523.700000 416.320000 524.180000 ;
        RECT 415.120000 518.260000 416.320000 518.740000 ;
        RECT 415.120000 512.820000 416.320000 513.300000 ;
        RECT 415.120000 507.380000 416.320000 507.860000 ;
        RECT 280.120000 529.140000 281.320000 529.620000 ;
        RECT 280.120000 534.580000 281.320000 535.060000 ;
        RECT 280.120000 540.020000 281.320000 540.500000 ;
        RECT 280.120000 561.780000 281.320000 562.260000 ;
        RECT 280.120000 556.340000 281.320000 556.820000 ;
        RECT 280.120000 550.900000 281.320000 551.380000 ;
        RECT 280.120000 545.460000 281.320000 545.940000 ;
        RECT 325.120000 529.140000 326.320000 529.620000 ;
        RECT 325.120000 534.580000 326.320000 535.060000 ;
        RECT 325.120000 540.020000 326.320000 540.500000 ;
        RECT 325.120000 561.780000 326.320000 562.260000 ;
        RECT 325.120000 556.340000 326.320000 556.820000 ;
        RECT 325.120000 550.900000 326.320000 551.380000 ;
        RECT 325.120000 545.460000 326.320000 545.940000 ;
        RECT 280.120000 567.220000 281.320000 567.700000 ;
        RECT 280.120000 572.660000 281.320000 573.140000 ;
        RECT 280.120000 578.100000 281.320000 578.580000 ;
        RECT 280.120000 583.540000 281.320000 584.020000 ;
        RECT 280.120000 588.980000 281.320000 589.460000 ;
        RECT 325.120000 567.220000 326.320000 567.700000 ;
        RECT 325.120000 572.660000 326.320000 573.140000 ;
        RECT 325.120000 578.100000 326.320000 578.580000 ;
        RECT 325.120000 583.540000 326.320000 584.020000 ;
        RECT 325.120000 588.980000 326.320000 589.460000 ;
        RECT 370.120000 529.140000 371.320000 529.620000 ;
        RECT 370.120000 534.580000 371.320000 535.060000 ;
        RECT 370.120000 540.020000 371.320000 540.500000 ;
        RECT 370.120000 561.780000 371.320000 562.260000 ;
        RECT 370.120000 556.340000 371.320000 556.820000 ;
        RECT 370.120000 550.900000 371.320000 551.380000 ;
        RECT 370.120000 545.460000 371.320000 545.940000 ;
        RECT 415.120000 529.140000 416.320000 529.620000 ;
        RECT 415.120000 534.580000 416.320000 535.060000 ;
        RECT 415.120000 540.020000 416.320000 540.500000 ;
        RECT 415.120000 561.780000 416.320000 562.260000 ;
        RECT 415.120000 556.340000 416.320000 556.820000 ;
        RECT 415.120000 550.900000 416.320000 551.380000 ;
        RECT 415.120000 545.460000 416.320000 545.940000 ;
        RECT 370.120000 567.220000 371.320000 567.700000 ;
        RECT 370.120000 572.660000 371.320000 573.140000 ;
        RECT 370.120000 578.100000 371.320000 578.580000 ;
        RECT 370.120000 583.540000 371.320000 584.020000 ;
        RECT 370.120000 588.980000 371.320000 589.460000 ;
        RECT 415.120000 567.220000 416.320000 567.700000 ;
        RECT 415.120000 572.660000 416.320000 573.140000 ;
        RECT 415.120000 578.100000 416.320000 578.580000 ;
        RECT 415.120000 583.540000 416.320000 584.020000 ;
        RECT 415.120000 588.980000 416.320000 589.460000 ;
        RECT 460.120000 485.620000 461.320000 486.100000 ;
        RECT 460.120000 480.180000 461.320000 480.660000 ;
        RECT 460.120000 474.740000 461.320000 475.220000 ;
        RECT 460.120000 469.300000 461.320000 469.780000 ;
        RECT 460.120000 452.980000 461.320000 453.460000 ;
        RECT 460.120000 458.420000 461.320000 458.900000 ;
        RECT 460.120000 463.860000 461.320000 464.340000 ;
        RECT 460.120000 523.700000 461.320000 524.180000 ;
        RECT 460.120000 518.260000 461.320000 518.740000 ;
        RECT 460.120000 512.820000 461.320000 513.300000 ;
        RECT 460.120000 507.380000 461.320000 507.860000 ;
        RECT 460.120000 491.060000 461.320000 491.540000 ;
        RECT 460.120000 496.500000 461.320000 496.980000 ;
        RECT 460.120000 501.940000 461.320000 502.420000 ;
        RECT 505.120000 463.860000 506.320000 464.340000 ;
        RECT 505.120000 458.420000 506.320000 458.900000 ;
        RECT 505.120000 452.980000 506.320000 453.460000 ;
        RECT 505.120000 485.620000 506.320000 486.100000 ;
        RECT 505.120000 480.180000 506.320000 480.660000 ;
        RECT 505.120000 474.740000 506.320000 475.220000 ;
        RECT 505.120000 469.300000 506.320000 469.780000 ;
        RECT 545.600000 463.860000 546.800000 464.340000 ;
        RECT 545.600000 458.420000 546.800000 458.900000 ;
        RECT 545.600000 452.980000 546.800000 453.460000 ;
        RECT 545.600000 485.620000 546.800000 486.100000 ;
        RECT 545.600000 480.180000 546.800000 480.660000 ;
        RECT 545.600000 474.740000 546.800000 475.220000 ;
        RECT 545.600000 469.300000 546.800000 469.780000 ;
        RECT 505.120000 501.940000 506.320000 502.420000 ;
        RECT 505.120000 496.500000 506.320000 496.980000 ;
        RECT 505.120000 491.060000 506.320000 491.540000 ;
        RECT 505.120000 523.700000 506.320000 524.180000 ;
        RECT 505.120000 518.260000 506.320000 518.740000 ;
        RECT 505.120000 512.820000 506.320000 513.300000 ;
        RECT 505.120000 507.380000 506.320000 507.860000 ;
        RECT 545.600000 501.940000 546.800000 502.420000 ;
        RECT 545.600000 496.500000 546.800000 496.980000 ;
        RECT 545.600000 491.060000 546.800000 491.540000 ;
        RECT 545.600000 523.700000 546.800000 524.180000 ;
        RECT 545.600000 518.260000 546.800000 518.740000 ;
        RECT 545.600000 512.820000 546.800000 513.300000 ;
        RECT 545.600000 507.380000 546.800000 507.860000 ;
        RECT 460.120000 561.780000 461.320000 562.260000 ;
        RECT 460.120000 556.340000 461.320000 556.820000 ;
        RECT 460.120000 550.900000 461.320000 551.380000 ;
        RECT 460.120000 545.460000 461.320000 545.940000 ;
        RECT 460.120000 529.140000 461.320000 529.620000 ;
        RECT 460.120000 534.580000 461.320000 535.060000 ;
        RECT 460.120000 540.020000 461.320000 540.500000 ;
        RECT 460.120000 567.220000 461.320000 567.700000 ;
        RECT 460.120000 572.660000 461.320000 573.140000 ;
        RECT 460.120000 578.100000 461.320000 578.580000 ;
        RECT 460.120000 583.540000 461.320000 584.020000 ;
        RECT 460.120000 588.980000 461.320000 589.460000 ;
        RECT 505.120000 540.020000 506.320000 540.500000 ;
        RECT 505.120000 534.580000 506.320000 535.060000 ;
        RECT 505.120000 529.140000 506.320000 529.620000 ;
        RECT 505.120000 561.780000 506.320000 562.260000 ;
        RECT 505.120000 556.340000 506.320000 556.820000 ;
        RECT 505.120000 550.900000 506.320000 551.380000 ;
        RECT 505.120000 545.460000 506.320000 545.940000 ;
        RECT 545.600000 540.020000 546.800000 540.500000 ;
        RECT 545.600000 534.580000 546.800000 535.060000 ;
        RECT 545.600000 529.140000 546.800000 529.620000 ;
        RECT 545.600000 561.780000 546.800000 562.260000 ;
        RECT 545.600000 556.340000 546.800000 556.820000 ;
        RECT 545.600000 550.900000 546.800000 551.380000 ;
        RECT 545.600000 545.460000 546.800000 545.940000 ;
        RECT 505.120000 578.100000 506.320000 578.580000 ;
        RECT 505.120000 572.660000 506.320000 573.140000 ;
        RECT 505.120000 567.220000 506.320000 567.700000 ;
        RECT 505.120000 583.540000 506.320000 584.020000 ;
        RECT 505.120000 588.980000 506.320000 589.460000 ;
        RECT 545.600000 578.100000 546.800000 578.580000 ;
        RECT 545.600000 567.220000 546.800000 567.700000 ;
        RECT 545.600000 572.660000 546.800000 573.140000 ;
        RECT 545.600000 588.980000 546.800000 589.460000 ;
        RECT 545.600000 583.540000 546.800000 584.020000 ;
      LAYER met4 ;
        RECT 505.120000 3.230000 506.320000 596.190000 ;
        RECT 460.120000 3.230000 461.320000 596.190000 ;
        RECT 415.120000 3.230000 416.320000 596.190000 ;
        RECT 370.120000 3.230000 371.320000 596.190000 ;
        RECT 325.120000 3.230000 326.320000 596.190000 ;
        RECT 280.120000 3.230000 281.320000 596.190000 ;
        RECT 235.120000 3.230000 236.320000 596.190000 ;
        RECT 190.120000 3.230000 191.320000 596.190000 ;
        RECT 145.120000 3.230000 146.320000 596.190000 ;
        RECT 100.120000 3.230000 101.320000 596.190000 ;
        RECT 55.120000 3.230000 56.320000 596.190000 ;
        RECT 10.120000 3.230000 11.320000 596.190000 ;
        RECT 545.600000 0.000000 546.800000 599.760000 ;
        RECT 3.360000 0.000000 4.560000 599.760000 ;
        RECT 9.955000 17.780000 11.320000 18.260000 ;
        RECT 9.955000 12.340000 11.320000 12.820000 ;
        RECT 9.955000 23.220000 11.320000 23.700000 ;
        RECT 9.955000 34.100000 11.320000 34.580000 ;
        RECT 9.955000 28.660000 11.320000 29.140000 ;
        RECT 9.955000 55.860000 11.320000 56.340000 ;
        RECT 9.955000 44.980000 11.320000 45.460000 ;
        RECT 9.955000 39.540000 11.320000 40.020000 ;
        RECT 9.955000 50.420000 11.320000 50.900000 ;
        RECT 9.955000 61.300000 11.320000 61.780000 ;
        RECT 9.955000 66.740000 11.320000 67.220000 ;
        RECT 9.955000 72.180000 11.320000 72.660000 ;
        RECT 9.955000 83.060000 11.320000 83.540000 ;
        RECT 9.955000 77.620000 11.320000 78.100000 ;
        RECT 9.955000 88.500000 11.320000 88.980000 ;
        RECT 9.955000 99.380000 11.320000 99.860000 ;
        RECT 9.955000 93.940000 11.320000 94.420000 ;
        RECT 9.955000 110.260000 11.320000 110.740000 ;
        RECT 9.955000 104.820000 11.320000 105.300000 ;
        RECT 9.955000 115.700000 11.320000 116.180000 ;
        RECT 9.955000 121.140000 11.320000 121.620000 ;
        RECT 9.955000 126.580000 11.320000 127.060000 ;
        RECT 9.955000 137.460000 11.320000 137.940000 ;
        RECT 9.955000 132.020000 11.320000 132.500000 ;
        RECT 9.955000 148.340000 11.320000 148.820000 ;
        RECT 9.955000 142.900000 11.320000 143.380000 ;
        RECT 9.955000 224.500000 11.320000 224.980000 ;
        RECT 9.955000 159.220000 11.320000 159.700000 ;
        RECT 9.955000 153.780000 11.320000 154.260000 ;
        RECT 9.955000 164.660000 11.320000 165.140000 ;
        RECT 9.955000 175.540000 11.320000 176.020000 ;
        RECT 9.955000 170.100000 11.320000 170.580000 ;
        RECT 9.955000 186.420000 11.320000 186.900000 ;
        RECT 9.955000 180.980000 11.320000 181.460000 ;
        RECT 9.955000 191.860000 11.320000 192.340000 ;
        RECT 9.955000 202.740000 11.320000 203.220000 ;
        RECT 9.955000 197.300000 11.320000 197.780000 ;
        RECT 9.955000 213.620000 11.320000 214.100000 ;
        RECT 9.955000 208.180000 11.320000 208.660000 ;
        RECT 9.955000 219.060000 11.320000 219.540000 ;
        RECT 9.955000 229.940000 11.320000 230.420000 ;
        RECT 9.955000 235.380000 11.320000 235.860000 ;
        RECT 9.955000 240.820000 11.320000 241.300000 ;
        RECT 9.955000 251.700000 11.320000 252.180000 ;
        RECT 9.955000 246.260000 11.320000 246.740000 ;
        RECT 9.955000 257.140000 11.320000 257.620000 ;
        RECT 9.955000 268.020000 11.320000 268.500000 ;
        RECT 9.955000 262.580000 11.320000 263.060000 ;
        RECT 9.955000 278.900000 11.320000 279.380000 ;
        RECT 9.955000 273.460000 11.320000 273.940000 ;
        RECT 9.955000 284.340000 11.320000 284.820000 ;
        RECT 9.955000 289.780000 11.320000 290.260000 ;
        RECT 9.955000 295.220000 11.320000 295.700000 ;
        RECT 9.955000 306.100000 11.320000 306.580000 ;
        RECT 9.955000 300.660000 11.320000 301.140000 ;
        RECT 9.955000 316.980000 11.320000 317.460000 ;
        RECT 9.955000 311.540000 11.320000 312.020000 ;
        RECT 9.955000 327.860000 11.320000 328.340000 ;
        RECT 9.955000 322.420000 11.320000 322.900000 ;
        RECT 9.955000 333.300000 11.320000 333.780000 ;
        RECT 9.955000 344.180000 11.320000 344.660000 ;
        RECT 9.955000 338.740000 11.320000 339.220000 ;
        RECT 9.955000 355.060000 11.320000 355.540000 ;
        RECT 9.955000 349.620000 11.320000 350.100000 ;
        RECT 9.955000 360.500000 11.320000 360.980000 ;
        RECT 9.955000 371.380000 11.320000 371.860000 ;
        RECT 9.955000 365.940000 11.320000 366.420000 ;
        RECT 9.955000 393.140000 11.320000 393.620000 ;
        RECT 9.955000 382.260000 11.320000 382.740000 ;
        RECT 9.955000 376.820000 11.320000 377.300000 ;
        RECT 9.955000 387.700000 11.320000 388.180000 ;
        RECT 9.955000 398.580000 11.320000 399.060000 ;
        RECT 9.955000 404.020000 11.320000 404.500000 ;
        RECT 9.955000 409.460000 11.320000 409.940000 ;
        RECT 9.955000 420.340000 11.320000 420.820000 ;
        RECT 9.955000 414.900000 11.320000 415.380000 ;
        RECT 9.955000 425.780000 11.320000 426.260000 ;
        RECT 9.955000 436.660000 11.320000 437.140000 ;
        RECT 9.955000 431.220000 11.320000 431.700000 ;
        RECT 9.955000 447.540000 11.320000 448.020000 ;
        RECT 9.955000 442.100000 11.320000 442.580000 ;
        RECT 9.955000 452.980000 11.320000 453.460000 ;
        RECT 9.955000 458.420000 11.320000 458.900000 ;
        RECT 9.955000 463.860000 11.320000 464.340000 ;
        RECT 9.955000 474.740000 11.320000 475.220000 ;
        RECT 9.955000 469.300000 11.320000 469.780000 ;
        RECT 9.955000 485.620000 11.320000 486.100000 ;
        RECT 9.955000 480.180000 11.320000 480.660000 ;
        RECT 9.955000 496.500000 11.320000 496.980000 ;
        RECT 9.955000 491.060000 11.320000 491.540000 ;
        RECT 9.955000 501.940000 11.320000 502.420000 ;
        RECT 9.955000 512.820000 11.320000 513.300000 ;
        RECT 9.955000 507.380000 11.320000 507.860000 ;
        RECT 9.955000 523.700000 11.320000 524.180000 ;
        RECT 9.955000 518.260000 11.320000 518.740000 ;
        RECT 9.955000 529.140000 11.320000 529.620000 ;
        RECT 9.955000 540.020000 11.320000 540.500000 ;
        RECT 9.955000 534.580000 11.320000 535.060000 ;
        RECT 9.955000 550.900000 11.320000 551.380000 ;
        RECT 9.955000 545.460000 11.320000 545.940000 ;
        RECT 9.955000 561.780000 11.320000 562.260000 ;
        RECT 9.955000 556.340000 11.320000 556.820000 ;
        RECT 9.955000 567.220000 11.320000 567.700000 ;
        RECT 9.955000 572.660000 11.320000 573.140000 ;
        RECT 9.955000 578.100000 11.320000 578.580000 ;
        RECT 9.955000 588.980000 11.320000 589.460000 ;
        RECT 9.955000 583.540000 11.320000 584.020000 ;
    END
# end of P/G power stripe data as pin

  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 550.160000 599.760000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 550.160000 599.760000 ;
    LAYER met2 ;
      RECT 0.000000 1.040000 550.160000 599.760000 ;
      RECT 539.680000 0.000000 550.160000 1.040000 ;
      RECT 538.760000 0.000000 539.020000 1.040000 ;
      RECT 537.380000 0.000000 538.100000 1.040000 ;
      RECT 536.000000 0.000000 536.720000 1.040000 ;
      RECT 534.620000 0.000000 535.340000 1.040000 ;
      RECT 533.700000 0.000000 533.960000 1.040000 ;
      RECT 532.320000 0.000000 533.040000 1.040000 ;
      RECT 530.940000 0.000000 531.660000 1.040000 ;
      RECT 529.560000 0.000000 530.280000 1.040000 ;
      RECT 528.180000 0.000000 528.900000 1.040000 ;
      RECT 527.260000 0.000000 527.520000 1.040000 ;
      RECT 525.880000 0.000000 526.600000 1.040000 ;
      RECT 524.500000 0.000000 525.220000 1.040000 ;
      RECT 523.120000 0.000000 523.840000 1.040000 ;
      RECT 522.200000 0.000000 522.460000 1.040000 ;
      RECT 520.820000 0.000000 521.540000 1.040000 ;
      RECT 519.440000 0.000000 520.160000 1.040000 ;
      RECT 518.060000 0.000000 518.780000 1.040000 ;
      RECT 516.680000 0.000000 517.400000 1.040000 ;
      RECT 515.760000 0.000000 516.020000 1.040000 ;
      RECT 514.380000 0.000000 515.100000 1.040000 ;
      RECT 513.000000 0.000000 513.720000 1.040000 ;
      RECT 511.620000 0.000000 512.340000 1.040000 ;
      RECT 510.700000 0.000000 510.960000 1.040000 ;
      RECT 509.320000 0.000000 510.040000 1.040000 ;
      RECT 507.940000 0.000000 508.660000 1.040000 ;
      RECT 506.560000 0.000000 507.280000 1.040000 ;
      RECT 505.180000 0.000000 505.900000 1.040000 ;
      RECT 504.260000 0.000000 504.520000 1.040000 ;
      RECT 502.880000 0.000000 503.600000 1.040000 ;
      RECT 501.500000 0.000000 502.220000 1.040000 ;
      RECT 500.120000 0.000000 500.840000 1.040000 ;
      RECT 499.200000 0.000000 499.460000 1.040000 ;
      RECT 497.820000 0.000000 498.540000 1.040000 ;
      RECT 496.440000 0.000000 497.160000 1.040000 ;
      RECT 495.060000 0.000000 495.780000 1.040000 ;
      RECT 493.680000 0.000000 494.400000 1.040000 ;
      RECT 492.760000 0.000000 493.020000 1.040000 ;
      RECT 491.380000 0.000000 492.100000 1.040000 ;
      RECT 490.000000 0.000000 490.720000 1.040000 ;
      RECT 488.620000 0.000000 489.340000 1.040000 ;
      RECT 487.700000 0.000000 487.960000 1.040000 ;
      RECT 486.320000 0.000000 487.040000 1.040000 ;
      RECT 484.940000 0.000000 485.660000 1.040000 ;
      RECT 483.560000 0.000000 484.280000 1.040000 ;
      RECT 482.180000 0.000000 482.900000 1.040000 ;
      RECT 481.260000 0.000000 481.520000 1.040000 ;
      RECT 479.880000 0.000000 480.600000 1.040000 ;
      RECT 478.500000 0.000000 479.220000 1.040000 ;
      RECT 477.120000 0.000000 477.840000 1.040000 ;
      RECT 475.740000 0.000000 476.460000 1.040000 ;
      RECT 474.820000 0.000000 475.080000 1.040000 ;
      RECT 473.440000 0.000000 474.160000 1.040000 ;
      RECT 472.060000 0.000000 472.780000 1.040000 ;
      RECT 470.680000 0.000000 471.400000 1.040000 ;
      RECT 469.760000 0.000000 470.020000 1.040000 ;
      RECT 468.380000 0.000000 469.100000 1.040000 ;
      RECT 467.000000 0.000000 467.720000 1.040000 ;
      RECT 465.620000 0.000000 466.340000 1.040000 ;
      RECT 464.240000 0.000000 464.960000 1.040000 ;
      RECT 463.320000 0.000000 463.580000 1.040000 ;
      RECT 461.940000 0.000000 462.660000 1.040000 ;
      RECT 460.560000 0.000000 461.280000 1.040000 ;
      RECT 459.180000 0.000000 459.900000 1.040000 ;
      RECT 458.260000 0.000000 458.520000 1.040000 ;
      RECT 456.880000 0.000000 457.600000 1.040000 ;
      RECT 455.500000 0.000000 456.220000 1.040000 ;
      RECT 454.120000 0.000000 454.840000 1.040000 ;
      RECT 452.740000 0.000000 453.460000 1.040000 ;
      RECT 451.820000 0.000000 452.080000 1.040000 ;
      RECT 450.440000 0.000000 451.160000 1.040000 ;
      RECT 449.060000 0.000000 449.780000 1.040000 ;
      RECT 447.680000 0.000000 448.400000 1.040000 ;
      RECT 446.760000 0.000000 447.020000 1.040000 ;
      RECT 445.380000 0.000000 446.100000 1.040000 ;
      RECT 444.000000 0.000000 444.720000 1.040000 ;
      RECT 442.620000 0.000000 443.340000 1.040000 ;
      RECT 441.240000 0.000000 441.960000 1.040000 ;
      RECT 440.320000 0.000000 440.580000 1.040000 ;
      RECT 438.940000 0.000000 439.660000 1.040000 ;
      RECT 437.560000 0.000000 438.280000 1.040000 ;
      RECT 436.180000 0.000000 436.900000 1.040000 ;
      RECT 435.260000 0.000000 435.520000 1.040000 ;
      RECT 433.880000 0.000000 434.600000 1.040000 ;
      RECT 432.500000 0.000000 433.220000 1.040000 ;
      RECT 431.120000 0.000000 431.840000 1.040000 ;
      RECT 429.740000 0.000000 430.460000 1.040000 ;
      RECT 428.820000 0.000000 429.080000 1.040000 ;
      RECT 427.440000 0.000000 428.160000 1.040000 ;
      RECT 426.060000 0.000000 426.780000 1.040000 ;
      RECT 424.680000 0.000000 425.400000 1.040000 ;
      RECT 423.760000 0.000000 424.020000 1.040000 ;
      RECT 422.380000 0.000000 423.100000 1.040000 ;
      RECT 421.000000 0.000000 421.720000 1.040000 ;
      RECT 419.620000 0.000000 420.340000 1.040000 ;
      RECT 418.240000 0.000000 418.960000 1.040000 ;
      RECT 417.320000 0.000000 417.580000 1.040000 ;
      RECT 415.940000 0.000000 416.660000 1.040000 ;
      RECT 414.560000 0.000000 415.280000 1.040000 ;
      RECT 413.180000 0.000000 413.900000 1.040000 ;
      RECT 411.800000 0.000000 412.520000 1.040000 ;
      RECT 410.880000 0.000000 411.140000 1.040000 ;
      RECT 409.500000 0.000000 410.220000 1.040000 ;
      RECT 408.120000 0.000000 408.840000 1.040000 ;
      RECT 406.740000 0.000000 407.460000 1.040000 ;
      RECT 405.820000 0.000000 406.080000 1.040000 ;
      RECT 404.440000 0.000000 405.160000 1.040000 ;
      RECT 403.060000 0.000000 403.780000 1.040000 ;
      RECT 401.680000 0.000000 402.400000 1.040000 ;
      RECT 400.300000 0.000000 401.020000 1.040000 ;
      RECT 399.380000 0.000000 399.640000 1.040000 ;
      RECT 398.000000 0.000000 398.720000 1.040000 ;
      RECT 396.620000 0.000000 397.340000 1.040000 ;
      RECT 395.240000 0.000000 395.960000 1.040000 ;
      RECT 394.320000 0.000000 394.580000 1.040000 ;
      RECT 392.940000 0.000000 393.660000 1.040000 ;
      RECT 391.560000 0.000000 392.280000 1.040000 ;
      RECT 390.180000 0.000000 390.900000 1.040000 ;
      RECT 388.800000 0.000000 389.520000 1.040000 ;
      RECT 387.880000 0.000000 388.140000 1.040000 ;
      RECT 386.500000 0.000000 387.220000 1.040000 ;
      RECT 385.120000 0.000000 385.840000 1.040000 ;
      RECT 383.740000 0.000000 384.460000 1.040000 ;
      RECT 382.820000 0.000000 383.080000 1.040000 ;
      RECT 381.440000 0.000000 382.160000 1.040000 ;
      RECT 380.060000 0.000000 380.780000 1.040000 ;
      RECT 378.680000 0.000000 379.400000 1.040000 ;
      RECT 377.300000 0.000000 378.020000 1.040000 ;
      RECT 376.380000 0.000000 376.640000 1.040000 ;
      RECT 375.000000 0.000000 375.720000 1.040000 ;
      RECT 373.620000 0.000000 374.340000 1.040000 ;
      RECT 372.240000 0.000000 372.960000 1.040000 ;
      RECT 371.320000 0.000000 371.580000 1.040000 ;
      RECT 369.940000 0.000000 370.660000 1.040000 ;
      RECT 368.560000 0.000000 369.280000 1.040000 ;
      RECT 367.180000 0.000000 367.900000 1.040000 ;
      RECT 365.800000 0.000000 366.520000 1.040000 ;
      RECT 364.880000 0.000000 365.140000 1.040000 ;
      RECT 363.500000 0.000000 364.220000 1.040000 ;
      RECT 362.120000 0.000000 362.840000 1.040000 ;
      RECT 360.740000 0.000000 361.460000 1.040000 ;
      RECT 359.360000 0.000000 360.080000 1.040000 ;
      RECT 358.440000 0.000000 358.700000 1.040000 ;
      RECT 357.060000 0.000000 357.780000 1.040000 ;
      RECT 355.680000 0.000000 356.400000 1.040000 ;
      RECT 354.300000 0.000000 355.020000 1.040000 ;
      RECT 353.380000 0.000000 353.640000 1.040000 ;
      RECT 352.000000 0.000000 352.720000 1.040000 ;
      RECT 350.620000 0.000000 351.340000 1.040000 ;
      RECT 349.240000 0.000000 349.960000 1.040000 ;
      RECT 347.860000 0.000000 348.580000 1.040000 ;
      RECT 346.940000 0.000000 347.200000 1.040000 ;
      RECT 345.560000 0.000000 346.280000 1.040000 ;
      RECT 344.180000 0.000000 344.900000 1.040000 ;
      RECT 342.800000 0.000000 343.520000 1.040000 ;
      RECT 341.880000 0.000000 342.140000 1.040000 ;
      RECT 340.500000 0.000000 341.220000 1.040000 ;
      RECT 339.120000 0.000000 339.840000 1.040000 ;
      RECT 337.740000 0.000000 338.460000 1.040000 ;
      RECT 336.360000 0.000000 337.080000 1.040000 ;
      RECT 335.440000 0.000000 335.700000 1.040000 ;
      RECT 334.060000 0.000000 334.780000 1.040000 ;
      RECT 332.680000 0.000000 333.400000 1.040000 ;
      RECT 331.300000 0.000000 332.020000 1.040000 ;
      RECT 330.380000 0.000000 330.640000 1.040000 ;
      RECT 329.000000 0.000000 329.720000 1.040000 ;
      RECT 327.620000 0.000000 328.340000 1.040000 ;
      RECT 326.240000 0.000000 326.960000 1.040000 ;
      RECT 324.860000 0.000000 325.580000 1.040000 ;
      RECT 323.940000 0.000000 324.200000 1.040000 ;
      RECT 322.560000 0.000000 323.280000 1.040000 ;
      RECT 321.180000 0.000000 321.900000 1.040000 ;
      RECT 319.800000 0.000000 320.520000 1.040000 ;
      RECT 318.880000 0.000000 319.140000 1.040000 ;
      RECT 317.500000 0.000000 318.220000 1.040000 ;
      RECT 316.120000 0.000000 316.840000 1.040000 ;
      RECT 314.740000 0.000000 315.460000 1.040000 ;
      RECT 313.360000 0.000000 314.080000 1.040000 ;
      RECT 312.440000 0.000000 312.700000 1.040000 ;
      RECT 311.060000 0.000000 311.780000 1.040000 ;
      RECT 309.680000 0.000000 310.400000 1.040000 ;
      RECT 308.300000 0.000000 309.020000 1.040000 ;
      RECT 307.380000 0.000000 307.640000 1.040000 ;
      RECT 306.000000 0.000000 306.720000 1.040000 ;
      RECT 304.620000 0.000000 305.340000 1.040000 ;
      RECT 303.240000 0.000000 303.960000 1.040000 ;
      RECT 301.860000 0.000000 302.580000 1.040000 ;
      RECT 300.940000 0.000000 301.200000 1.040000 ;
      RECT 299.560000 0.000000 300.280000 1.040000 ;
      RECT 298.180000 0.000000 298.900000 1.040000 ;
      RECT 296.800000 0.000000 297.520000 1.040000 ;
      RECT 295.420000 0.000000 296.140000 1.040000 ;
      RECT 294.500000 0.000000 294.760000 1.040000 ;
      RECT 293.120000 0.000000 293.840000 1.040000 ;
      RECT 291.740000 0.000000 292.460000 1.040000 ;
      RECT 290.360000 0.000000 291.080000 1.040000 ;
      RECT 289.440000 0.000000 289.700000 1.040000 ;
      RECT 288.060000 0.000000 288.780000 1.040000 ;
      RECT 286.680000 0.000000 287.400000 1.040000 ;
      RECT 285.300000 0.000000 286.020000 1.040000 ;
      RECT 283.920000 0.000000 284.640000 1.040000 ;
      RECT 283.000000 0.000000 283.260000 1.040000 ;
      RECT 281.620000 0.000000 282.340000 1.040000 ;
      RECT 280.240000 0.000000 280.960000 1.040000 ;
      RECT 278.860000 0.000000 279.580000 1.040000 ;
      RECT 277.940000 0.000000 278.200000 1.040000 ;
      RECT 276.560000 0.000000 277.280000 1.040000 ;
      RECT 275.180000 0.000000 275.900000 1.040000 ;
      RECT 273.800000 0.000000 274.520000 1.040000 ;
      RECT 272.420000 0.000000 273.140000 1.040000 ;
      RECT 271.500000 0.000000 271.760000 1.040000 ;
      RECT 270.120000 0.000000 270.840000 1.040000 ;
      RECT 268.740000 0.000000 269.460000 1.040000 ;
      RECT 267.360000 0.000000 268.080000 1.040000 ;
      RECT 266.440000 0.000000 266.700000 1.040000 ;
      RECT 265.060000 0.000000 265.780000 1.040000 ;
      RECT 263.680000 0.000000 264.400000 1.040000 ;
      RECT 262.300000 0.000000 263.020000 1.040000 ;
      RECT 260.920000 0.000000 261.640000 1.040000 ;
      RECT 260.000000 0.000000 260.260000 1.040000 ;
      RECT 258.620000 0.000000 259.340000 1.040000 ;
      RECT 257.240000 0.000000 257.960000 1.040000 ;
      RECT 255.860000 0.000000 256.580000 1.040000 ;
      RECT 254.940000 0.000000 255.200000 1.040000 ;
      RECT 253.560000 0.000000 254.280000 1.040000 ;
      RECT 252.180000 0.000000 252.900000 1.040000 ;
      RECT 250.800000 0.000000 251.520000 1.040000 ;
      RECT 249.420000 0.000000 250.140000 1.040000 ;
      RECT 248.500000 0.000000 248.760000 1.040000 ;
      RECT 247.120000 0.000000 247.840000 1.040000 ;
      RECT 245.740000 0.000000 246.460000 1.040000 ;
      RECT 244.360000 0.000000 245.080000 1.040000 ;
      RECT 242.980000 0.000000 243.700000 1.040000 ;
      RECT 242.060000 0.000000 242.320000 1.040000 ;
      RECT 240.680000 0.000000 241.400000 1.040000 ;
      RECT 239.300000 0.000000 240.020000 1.040000 ;
      RECT 237.920000 0.000000 238.640000 1.040000 ;
      RECT 237.000000 0.000000 237.260000 1.040000 ;
      RECT 235.620000 0.000000 236.340000 1.040000 ;
      RECT 234.240000 0.000000 234.960000 1.040000 ;
      RECT 232.860000 0.000000 233.580000 1.040000 ;
      RECT 231.480000 0.000000 232.200000 1.040000 ;
      RECT 230.560000 0.000000 230.820000 1.040000 ;
      RECT 229.180000 0.000000 229.900000 1.040000 ;
      RECT 227.800000 0.000000 228.520000 1.040000 ;
      RECT 226.420000 0.000000 227.140000 1.040000 ;
      RECT 225.500000 0.000000 225.760000 1.040000 ;
      RECT 224.120000 0.000000 224.840000 1.040000 ;
      RECT 222.740000 0.000000 223.460000 1.040000 ;
      RECT 221.360000 0.000000 222.080000 1.040000 ;
      RECT 219.980000 0.000000 220.700000 1.040000 ;
      RECT 219.060000 0.000000 219.320000 1.040000 ;
      RECT 217.680000 0.000000 218.400000 1.040000 ;
      RECT 216.300000 0.000000 217.020000 1.040000 ;
      RECT 214.920000 0.000000 215.640000 1.040000 ;
      RECT 214.000000 0.000000 214.260000 1.040000 ;
      RECT 212.620000 0.000000 213.340000 1.040000 ;
      RECT 211.240000 0.000000 211.960000 1.040000 ;
      RECT 209.860000 0.000000 210.580000 1.040000 ;
      RECT 208.480000 0.000000 209.200000 1.040000 ;
      RECT 207.560000 0.000000 207.820000 1.040000 ;
      RECT 206.180000 0.000000 206.900000 1.040000 ;
      RECT 204.800000 0.000000 205.520000 1.040000 ;
      RECT 203.420000 0.000000 204.140000 1.040000 ;
      RECT 202.500000 0.000000 202.760000 1.040000 ;
      RECT 201.120000 0.000000 201.840000 1.040000 ;
      RECT 199.740000 0.000000 200.460000 1.040000 ;
      RECT 198.360000 0.000000 199.080000 1.040000 ;
      RECT 196.980000 0.000000 197.700000 1.040000 ;
      RECT 196.060000 0.000000 196.320000 1.040000 ;
      RECT 194.680000 0.000000 195.400000 1.040000 ;
      RECT 193.300000 0.000000 194.020000 1.040000 ;
      RECT 191.920000 0.000000 192.640000 1.040000 ;
      RECT 191.000000 0.000000 191.260000 1.040000 ;
      RECT 189.620000 0.000000 190.340000 1.040000 ;
      RECT 188.240000 0.000000 188.960000 1.040000 ;
      RECT 186.860000 0.000000 187.580000 1.040000 ;
      RECT 185.480000 0.000000 186.200000 1.040000 ;
      RECT 184.560000 0.000000 184.820000 1.040000 ;
      RECT 183.180000 0.000000 183.900000 1.040000 ;
      RECT 181.800000 0.000000 182.520000 1.040000 ;
      RECT 180.420000 0.000000 181.140000 1.040000 ;
      RECT 179.040000 0.000000 179.760000 1.040000 ;
      RECT 178.120000 0.000000 178.380000 1.040000 ;
      RECT 176.740000 0.000000 177.460000 1.040000 ;
      RECT 175.360000 0.000000 176.080000 1.040000 ;
      RECT 173.980000 0.000000 174.700000 1.040000 ;
      RECT 173.060000 0.000000 173.320000 1.040000 ;
      RECT 171.680000 0.000000 172.400000 1.040000 ;
      RECT 170.300000 0.000000 171.020000 1.040000 ;
      RECT 168.920000 0.000000 169.640000 1.040000 ;
      RECT 167.540000 0.000000 168.260000 1.040000 ;
      RECT 166.620000 0.000000 166.880000 1.040000 ;
      RECT 165.240000 0.000000 165.960000 1.040000 ;
      RECT 163.860000 0.000000 164.580000 1.040000 ;
      RECT 162.480000 0.000000 163.200000 1.040000 ;
      RECT 161.560000 0.000000 161.820000 1.040000 ;
      RECT 160.180000 0.000000 160.900000 1.040000 ;
      RECT 158.800000 0.000000 159.520000 1.040000 ;
      RECT 157.420000 0.000000 158.140000 1.040000 ;
      RECT 156.040000 0.000000 156.760000 1.040000 ;
      RECT 155.120000 0.000000 155.380000 1.040000 ;
      RECT 153.740000 0.000000 154.460000 1.040000 ;
      RECT 152.360000 0.000000 153.080000 1.040000 ;
      RECT 150.980000 0.000000 151.700000 1.040000 ;
      RECT 150.060000 0.000000 150.320000 1.040000 ;
      RECT 148.680000 0.000000 149.400000 1.040000 ;
      RECT 147.300000 0.000000 148.020000 1.040000 ;
      RECT 145.920000 0.000000 146.640000 1.040000 ;
      RECT 144.540000 0.000000 145.260000 1.040000 ;
      RECT 143.620000 0.000000 143.880000 1.040000 ;
      RECT 142.240000 0.000000 142.960000 1.040000 ;
      RECT 140.860000 0.000000 141.580000 1.040000 ;
      RECT 139.480000 0.000000 140.200000 1.040000 ;
      RECT 138.560000 0.000000 138.820000 1.040000 ;
      RECT 137.180000 0.000000 137.900000 1.040000 ;
      RECT 135.800000 0.000000 136.520000 1.040000 ;
      RECT 134.420000 0.000000 135.140000 1.040000 ;
      RECT 133.040000 0.000000 133.760000 1.040000 ;
      RECT 132.120000 0.000000 132.380000 1.040000 ;
      RECT 130.740000 0.000000 131.460000 1.040000 ;
      RECT 129.360000 0.000000 130.080000 1.040000 ;
      RECT 127.980000 0.000000 128.700000 1.040000 ;
      RECT 126.600000 0.000000 127.320000 1.040000 ;
      RECT 125.680000 0.000000 125.940000 1.040000 ;
      RECT 124.300000 0.000000 125.020000 1.040000 ;
      RECT 122.920000 0.000000 123.640000 1.040000 ;
      RECT 121.540000 0.000000 122.260000 1.040000 ;
      RECT 120.620000 0.000000 120.880000 1.040000 ;
      RECT 119.240000 0.000000 119.960000 1.040000 ;
      RECT 117.860000 0.000000 118.580000 1.040000 ;
      RECT 116.480000 0.000000 117.200000 1.040000 ;
      RECT 115.100000 0.000000 115.820000 1.040000 ;
      RECT 114.180000 0.000000 114.440000 1.040000 ;
      RECT 112.800000 0.000000 113.520000 1.040000 ;
      RECT 111.420000 0.000000 112.140000 1.040000 ;
      RECT 110.040000 0.000000 110.760000 1.040000 ;
      RECT 109.120000 0.000000 109.380000 1.040000 ;
      RECT 107.740000 0.000000 108.460000 1.040000 ;
      RECT 106.360000 0.000000 107.080000 1.040000 ;
      RECT 104.980000 0.000000 105.700000 1.040000 ;
      RECT 103.600000 0.000000 104.320000 1.040000 ;
      RECT 102.680000 0.000000 102.940000 1.040000 ;
      RECT 101.300000 0.000000 102.020000 1.040000 ;
      RECT 99.920000 0.000000 100.640000 1.040000 ;
      RECT 98.540000 0.000000 99.260000 1.040000 ;
      RECT 97.620000 0.000000 97.880000 1.040000 ;
      RECT 96.240000 0.000000 96.960000 1.040000 ;
      RECT 94.860000 0.000000 95.580000 1.040000 ;
      RECT 93.480000 0.000000 94.200000 1.040000 ;
      RECT 92.100000 0.000000 92.820000 1.040000 ;
      RECT 91.180000 0.000000 91.440000 1.040000 ;
      RECT 89.800000 0.000000 90.520000 1.040000 ;
      RECT 88.420000 0.000000 89.140000 1.040000 ;
      RECT 87.040000 0.000000 87.760000 1.040000 ;
      RECT 86.120000 0.000000 86.380000 1.040000 ;
      RECT 84.740000 0.000000 85.460000 1.040000 ;
      RECT 83.360000 0.000000 84.080000 1.040000 ;
      RECT 81.980000 0.000000 82.700000 1.040000 ;
      RECT 80.600000 0.000000 81.320000 1.040000 ;
      RECT 79.680000 0.000000 79.940000 1.040000 ;
      RECT 78.300000 0.000000 79.020000 1.040000 ;
      RECT 76.920000 0.000000 77.640000 1.040000 ;
      RECT 75.540000 0.000000 76.260000 1.040000 ;
      RECT 74.620000 0.000000 74.880000 1.040000 ;
      RECT 73.240000 0.000000 73.960000 1.040000 ;
      RECT 71.860000 0.000000 72.580000 1.040000 ;
      RECT 70.480000 0.000000 71.200000 1.040000 ;
      RECT 69.100000 0.000000 69.820000 1.040000 ;
      RECT 68.180000 0.000000 68.440000 1.040000 ;
      RECT 66.800000 0.000000 67.520000 1.040000 ;
      RECT 65.420000 0.000000 66.140000 1.040000 ;
      RECT 64.040000 0.000000 64.760000 1.040000 ;
      RECT 62.660000 0.000000 63.380000 1.040000 ;
      RECT 61.740000 0.000000 62.000000 1.040000 ;
      RECT 60.360000 0.000000 61.080000 1.040000 ;
      RECT 58.980000 0.000000 59.700000 1.040000 ;
      RECT 57.600000 0.000000 58.320000 1.040000 ;
      RECT 56.680000 0.000000 56.940000 1.040000 ;
      RECT 55.300000 0.000000 56.020000 1.040000 ;
      RECT 53.920000 0.000000 54.640000 1.040000 ;
      RECT 52.540000 0.000000 53.260000 1.040000 ;
      RECT 51.160000 0.000000 51.880000 1.040000 ;
      RECT 50.240000 0.000000 50.500000 1.040000 ;
      RECT 48.860000 0.000000 49.580000 1.040000 ;
      RECT 47.480000 0.000000 48.200000 1.040000 ;
      RECT 46.100000 0.000000 46.820000 1.040000 ;
      RECT 45.180000 0.000000 45.440000 1.040000 ;
      RECT 43.800000 0.000000 44.520000 1.040000 ;
      RECT 42.420000 0.000000 43.140000 1.040000 ;
      RECT 41.040000 0.000000 41.760000 1.040000 ;
      RECT 39.660000 0.000000 40.380000 1.040000 ;
      RECT 38.740000 0.000000 39.000000 1.040000 ;
      RECT 37.360000 0.000000 38.080000 1.040000 ;
      RECT 35.980000 0.000000 36.700000 1.040000 ;
      RECT 34.600000 0.000000 35.320000 1.040000 ;
      RECT 33.680000 0.000000 33.940000 1.040000 ;
      RECT 32.300000 0.000000 33.020000 1.040000 ;
      RECT 30.920000 0.000000 31.640000 1.040000 ;
      RECT 29.540000 0.000000 30.260000 1.040000 ;
      RECT 28.160000 0.000000 28.880000 1.040000 ;
      RECT 27.240000 0.000000 27.500000 1.040000 ;
      RECT 25.860000 0.000000 26.580000 1.040000 ;
      RECT 24.480000 0.000000 25.200000 1.040000 ;
      RECT 23.100000 0.000000 23.820000 1.040000 ;
      RECT 22.180000 0.000000 22.440000 1.040000 ;
      RECT 20.800000 0.000000 21.520000 1.040000 ;
      RECT 19.420000 0.000000 20.140000 1.040000 ;
      RECT 18.040000 0.000000 18.760000 1.040000 ;
      RECT 16.660000 0.000000 17.380000 1.040000 ;
      RECT 15.740000 0.000000 16.000000 1.040000 ;
      RECT 14.360000 0.000000 15.080000 1.040000 ;
      RECT 12.980000 0.000000 13.700000 1.040000 ;
      RECT 11.600000 0.000000 12.320000 1.040000 ;
      RECT 10.680000 0.000000 10.940000 1.040000 ;
      RECT 0.000000 0.000000 10.020000 1.040000 ;
    LAYER met3 ;
      RECT 0.000000 596.490000 550.160000 599.760000 ;
      RECT 0.000000 594.290000 550.160000 594.690000 ;
      RECT 0.000000 590.020000 550.160000 592.490000 ;
      RECT 0.000000 589.760000 548.960000 590.020000 ;
      RECT 547.100000 589.040000 548.960000 589.760000 ;
      RECT 547.100000 588.680000 550.160000 589.040000 ;
      RECT 506.620000 588.680000 545.300000 589.760000 ;
      RECT 461.620000 588.680000 504.820000 589.760000 ;
      RECT 416.620000 588.680000 459.820000 589.760000 ;
      RECT 371.620000 588.680000 414.820000 589.760000 ;
      RECT 326.620000 588.680000 369.820000 589.760000 ;
      RECT 281.620000 588.680000 324.820000 589.760000 ;
      RECT 236.620000 588.680000 279.820000 589.760000 ;
      RECT 191.620000 588.680000 234.820000 589.760000 ;
      RECT 146.620000 588.680000 189.820000 589.760000 ;
      RECT 101.620000 588.680000 144.820000 589.760000 ;
      RECT 56.620000 588.680000 99.820000 589.760000 ;
      RECT 11.620000 588.680000 54.820000 589.760000 ;
      RECT 4.860000 588.680000 9.655000 589.760000 ;
      RECT 0.000000 588.680000 3.060000 589.760000 ;
      RECT 0.000000 587.040000 550.160000 588.680000 ;
      RECT 544.900000 586.360000 550.160000 587.040000 ;
      RECT 544.900000 585.960000 548.960000 586.360000 ;
      RECT 508.620000 585.960000 543.100000 587.040000 ;
      RECT 463.620000 585.960000 506.820000 587.040000 ;
      RECT 418.620000 585.960000 461.820000 587.040000 ;
      RECT 373.620000 585.960000 416.820000 587.040000 ;
      RECT 328.620000 585.960000 371.820000 587.040000 ;
      RECT 283.620000 585.960000 326.820000 587.040000 ;
      RECT 238.620000 585.960000 281.820000 587.040000 ;
      RECT 193.620000 585.960000 236.820000 587.040000 ;
      RECT 148.620000 585.960000 191.820000 587.040000 ;
      RECT 103.620000 585.960000 146.820000 587.040000 ;
      RECT 58.620000 585.960000 101.820000 587.040000 ;
      RECT 13.620000 585.960000 56.820000 587.040000 ;
      RECT 7.060000 585.960000 11.820000 587.040000 ;
      RECT 0.000000 585.960000 5.260000 587.040000 ;
      RECT 0.000000 585.380000 548.960000 585.960000 ;
      RECT 0.000000 584.320000 550.160000 585.380000 ;
      RECT 547.100000 583.240000 550.160000 584.320000 ;
      RECT 506.620000 583.240000 545.300000 584.320000 ;
      RECT 461.620000 583.240000 504.820000 584.320000 ;
      RECT 416.620000 583.240000 459.820000 584.320000 ;
      RECT 371.620000 583.240000 414.820000 584.320000 ;
      RECT 326.620000 583.240000 369.820000 584.320000 ;
      RECT 281.620000 583.240000 324.820000 584.320000 ;
      RECT 236.620000 583.240000 279.820000 584.320000 ;
      RECT 191.620000 583.240000 234.820000 584.320000 ;
      RECT 146.620000 583.240000 189.820000 584.320000 ;
      RECT 101.620000 583.240000 144.820000 584.320000 ;
      RECT 56.620000 583.240000 99.820000 584.320000 ;
      RECT 11.620000 583.240000 54.820000 584.320000 ;
      RECT 4.860000 583.240000 9.655000 584.320000 ;
      RECT 0.000000 583.240000 3.060000 584.320000 ;
      RECT 0.000000 582.700000 550.160000 583.240000 ;
      RECT 0.000000 581.720000 548.960000 582.700000 ;
      RECT 0.000000 581.600000 550.160000 581.720000 ;
      RECT 544.900000 580.520000 550.160000 581.600000 ;
      RECT 508.620000 580.520000 543.100000 581.600000 ;
      RECT 463.620000 580.520000 506.820000 581.600000 ;
      RECT 418.620000 580.520000 461.820000 581.600000 ;
      RECT 373.620000 580.520000 416.820000 581.600000 ;
      RECT 328.620000 580.520000 371.820000 581.600000 ;
      RECT 283.620000 580.520000 326.820000 581.600000 ;
      RECT 238.620000 580.520000 281.820000 581.600000 ;
      RECT 193.620000 580.520000 236.820000 581.600000 ;
      RECT 148.620000 580.520000 191.820000 581.600000 ;
      RECT 103.620000 580.520000 146.820000 581.600000 ;
      RECT 58.620000 580.520000 101.820000 581.600000 ;
      RECT 13.620000 580.520000 56.820000 581.600000 ;
      RECT 7.060000 580.520000 11.820000 581.600000 ;
      RECT 0.000000 580.520000 5.260000 581.600000 ;
      RECT 0.000000 579.650000 550.160000 580.520000 ;
      RECT 0.000000 578.880000 548.960000 579.650000 ;
      RECT 547.100000 578.670000 548.960000 578.880000 ;
      RECT 547.100000 577.800000 550.160000 578.670000 ;
      RECT 506.620000 577.800000 545.300000 578.880000 ;
      RECT 461.620000 577.800000 504.820000 578.880000 ;
      RECT 416.620000 577.800000 459.820000 578.880000 ;
      RECT 371.620000 577.800000 414.820000 578.880000 ;
      RECT 326.620000 577.800000 369.820000 578.880000 ;
      RECT 281.620000 577.800000 324.820000 578.880000 ;
      RECT 236.620000 577.800000 279.820000 578.880000 ;
      RECT 191.620000 577.800000 234.820000 578.880000 ;
      RECT 146.620000 577.800000 189.820000 578.880000 ;
      RECT 101.620000 577.800000 144.820000 578.880000 ;
      RECT 56.620000 577.800000 99.820000 578.880000 ;
      RECT 11.620000 577.800000 54.820000 578.880000 ;
      RECT 4.860000 577.800000 9.655000 578.880000 ;
      RECT 0.000000 577.800000 3.060000 578.880000 ;
      RECT 0.000000 576.160000 550.160000 577.800000 ;
      RECT 544.900000 575.990000 550.160000 576.160000 ;
      RECT 544.900000 575.080000 548.960000 575.990000 ;
      RECT 508.620000 575.080000 543.100000 576.160000 ;
      RECT 463.620000 575.080000 506.820000 576.160000 ;
      RECT 418.620000 575.080000 461.820000 576.160000 ;
      RECT 373.620000 575.080000 416.820000 576.160000 ;
      RECT 328.620000 575.080000 371.820000 576.160000 ;
      RECT 283.620000 575.080000 326.820000 576.160000 ;
      RECT 238.620000 575.080000 281.820000 576.160000 ;
      RECT 193.620000 575.080000 236.820000 576.160000 ;
      RECT 148.620000 575.080000 191.820000 576.160000 ;
      RECT 103.620000 575.080000 146.820000 576.160000 ;
      RECT 58.620000 575.080000 101.820000 576.160000 ;
      RECT 13.620000 575.080000 56.820000 576.160000 ;
      RECT 7.060000 575.080000 11.820000 576.160000 ;
      RECT 0.000000 575.080000 5.260000 576.160000 ;
      RECT 0.000000 575.010000 548.960000 575.080000 ;
      RECT 0.000000 573.440000 550.160000 575.010000 ;
      RECT 547.100000 572.360000 550.160000 573.440000 ;
      RECT 506.620000 572.360000 545.300000 573.440000 ;
      RECT 461.620000 572.360000 504.820000 573.440000 ;
      RECT 416.620000 572.360000 459.820000 573.440000 ;
      RECT 371.620000 572.360000 414.820000 573.440000 ;
      RECT 326.620000 572.360000 369.820000 573.440000 ;
      RECT 281.620000 572.360000 324.820000 573.440000 ;
      RECT 236.620000 572.360000 279.820000 573.440000 ;
      RECT 191.620000 572.360000 234.820000 573.440000 ;
      RECT 146.620000 572.360000 189.820000 573.440000 ;
      RECT 101.620000 572.360000 144.820000 573.440000 ;
      RECT 56.620000 572.360000 99.820000 573.440000 ;
      RECT 11.620000 572.360000 54.820000 573.440000 ;
      RECT 4.860000 572.360000 9.655000 573.440000 ;
      RECT 0.000000 572.360000 3.060000 573.440000 ;
      RECT 0.000000 572.330000 550.160000 572.360000 ;
      RECT 0.000000 571.350000 548.960000 572.330000 ;
      RECT 0.000000 570.720000 550.160000 571.350000 ;
      RECT 544.900000 569.640000 550.160000 570.720000 ;
      RECT 508.620000 569.640000 543.100000 570.720000 ;
      RECT 463.620000 569.640000 506.820000 570.720000 ;
      RECT 418.620000 569.640000 461.820000 570.720000 ;
      RECT 373.620000 569.640000 416.820000 570.720000 ;
      RECT 328.620000 569.640000 371.820000 570.720000 ;
      RECT 283.620000 569.640000 326.820000 570.720000 ;
      RECT 238.620000 569.640000 281.820000 570.720000 ;
      RECT 193.620000 569.640000 236.820000 570.720000 ;
      RECT 148.620000 569.640000 191.820000 570.720000 ;
      RECT 103.620000 569.640000 146.820000 570.720000 ;
      RECT 58.620000 569.640000 101.820000 570.720000 ;
      RECT 13.620000 569.640000 56.820000 570.720000 ;
      RECT 7.060000 569.640000 11.820000 570.720000 ;
      RECT 0.000000 569.640000 5.260000 570.720000 ;
      RECT 0.000000 569.280000 550.160000 569.640000 ;
      RECT 0.000000 568.300000 548.960000 569.280000 ;
      RECT 0.000000 568.000000 550.160000 568.300000 ;
      RECT 547.100000 566.920000 550.160000 568.000000 ;
      RECT 506.620000 566.920000 545.300000 568.000000 ;
      RECT 461.620000 566.920000 504.820000 568.000000 ;
      RECT 416.620000 566.920000 459.820000 568.000000 ;
      RECT 371.620000 566.920000 414.820000 568.000000 ;
      RECT 326.620000 566.920000 369.820000 568.000000 ;
      RECT 281.620000 566.920000 324.820000 568.000000 ;
      RECT 236.620000 566.920000 279.820000 568.000000 ;
      RECT 191.620000 566.920000 234.820000 568.000000 ;
      RECT 146.620000 566.920000 189.820000 568.000000 ;
      RECT 101.620000 566.920000 144.820000 568.000000 ;
      RECT 56.620000 566.920000 99.820000 568.000000 ;
      RECT 11.620000 566.920000 54.820000 568.000000 ;
      RECT 4.860000 566.920000 9.655000 568.000000 ;
      RECT 0.000000 566.920000 3.060000 568.000000 ;
      RECT 0.000000 565.620000 550.160000 566.920000 ;
      RECT 0.000000 565.280000 548.960000 565.620000 ;
      RECT 544.900000 564.640000 548.960000 565.280000 ;
      RECT 544.900000 564.200000 550.160000 564.640000 ;
      RECT 508.620000 564.200000 543.100000 565.280000 ;
      RECT 463.620000 564.200000 506.820000 565.280000 ;
      RECT 418.620000 564.200000 461.820000 565.280000 ;
      RECT 373.620000 564.200000 416.820000 565.280000 ;
      RECT 328.620000 564.200000 371.820000 565.280000 ;
      RECT 283.620000 564.200000 326.820000 565.280000 ;
      RECT 238.620000 564.200000 281.820000 565.280000 ;
      RECT 193.620000 564.200000 236.820000 565.280000 ;
      RECT 148.620000 564.200000 191.820000 565.280000 ;
      RECT 103.620000 564.200000 146.820000 565.280000 ;
      RECT 58.620000 564.200000 101.820000 565.280000 ;
      RECT 13.620000 564.200000 56.820000 565.280000 ;
      RECT 7.060000 564.200000 11.820000 565.280000 ;
      RECT 0.000000 564.200000 5.260000 565.280000 ;
      RECT 0.000000 562.560000 550.160000 564.200000 ;
      RECT 547.100000 561.960000 550.160000 562.560000 ;
      RECT 547.100000 561.480000 548.960000 561.960000 ;
      RECT 506.620000 561.480000 545.300000 562.560000 ;
      RECT 461.620000 561.480000 504.820000 562.560000 ;
      RECT 416.620000 561.480000 459.820000 562.560000 ;
      RECT 371.620000 561.480000 414.820000 562.560000 ;
      RECT 326.620000 561.480000 369.820000 562.560000 ;
      RECT 281.620000 561.480000 324.820000 562.560000 ;
      RECT 236.620000 561.480000 279.820000 562.560000 ;
      RECT 191.620000 561.480000 234.820000 562.560000 ;
      RECT 146.620000 561.480000 189.820000 562.560000 ;
      RECT 101.620000 561.480000 144.820000 562.560000 ;
      RECT 56.620000 561.480000 99.820000 562.560000 ;
      RECT 11.620000 561.480000 54.820000 562.560000 ;
      RECT 4.860000 561.480000 9.655000 562.560000 ;
      RECT 0.000000 561.480000 3.060000 562.560000 ;
      RECT 0.000000 560.980000 548.960000 561.480000 ;
      RECT 0.000000 559.840000 550.160000 560.980000 ;
      RECT 544.900000 558.910000 550.160000 559.840000 ;
      RECT 544.900000 558.760000 548.960000 558.910000 ;
      RECT 508.620000 558.760000 543.100000 559.840000 ;
      RECT 463.620000 558.760000 506.820000 559.840000 ;
      RECT 418.620000 558.760000 461.820000 559.840000 ;
      RECT 373.620000 558.760000 416.820000 559.840000 ;
      RECT 328.620000 558.760000 371.820000 559.840000 ;
      RECT 283.620000 558.760000 326.820000 559.840000 ;
      RECT 238.620000 558.760000 281.820000 559.840000 ;
      RECT 193.620000 558.760000 236.820000 559.840000 ;
      RECT 148.620000 558.760000 191.820000 559.840000 ;
      RECT 103.620000 558.760000 146.820000 559.840000 ;
      RECT 58.620000 558.760000 101.820000 559.840000 ;
      RECT 13.620000 558.760000 56.820000 559.840000 ;
      RECT 7.060000 558.760000 11.820000 559.840000 ;
      RECT 0.000000 558.760000 5.260000 559.840000 ;
      RECT 0.000000 557.930000 548.960000 558.760000 ;
      RECT 0.000000 557.120000 550.160000 557.930000 ;
      RECT 547.100000 556.040000 550.160000 557.120000 ;
      RECT 506.620000 556.040000 545.300000 557.120000 ;
      RECT 461.620000 556.040000 504.820000 557.120000 ;
      RECT 416.620000 556.040000 459.820000 557.120000 ;
      RECT 371.620000 556.040000 414.820000 557.120000 ;
      RECT 326.620000 556.040000 369.820000 557.120000 ;
      RECT 281.620000 556.040000 324.820000 557.120000 ;
      RECT 236.620000 556.040000 279.820000 557.120000 ;
      RECT 191.620000 556.040000 234.820000 557.120000 ;
      RECT 146.620000 556.040000 189.820000 557.120000 ;
      RECT 101.620000 556.040000 144.820000 557.120000 ;
      RECT 56.620000 556.040000 99.820000 557.120000 ;
      RECT 11.620000 556.040000 54.820000 557.120000 ;
      RECT 4.860000 556.040000 9.655000 557.120000 ;
      RECT 0.000000 556.040000 3.060000 557.120000 ;
      RECT 0.000000 555.250000 550.160000 556.040000 ;
      RECT 0.000000 554.400000 548.960000 555.250000 ;
      RECT 544.900000 554.270000 548.960000 554.400000 ;
      RECT 544.900000 553.320000 550.160000 554.270000 ;
      RECT 508.620000 553.320000 543.100000 554.400000 ;
      RECT 463.620000 553.320000 506.820000 554.400000 ;
      RECT 418.620000 553.320000 461.820000 554.400000 ;
      RECT 373.620000 553.320000 416.820000 554.400000 ;
      RECT 328.620000 553.320000 371.820000 554.400000 ;
      RECT 283.620000 553.320000 326.820000 554.400000 ;
      RECT 238.620000 553.320000 281.820000 554.400000 ;
      RECT 193.620000 553.320000 236.820000 554.400000 ;
      RECT 148.620000 553.320000 191.820000 554.400000 ;
      RECT 103.620000 553.320000 146.820000 554.400000 ;
      RECT 58.620000 553.320000 101.820000 554.400000 ;
      RECT 13.620000 553.320000 56.820000 554.400000 ;
      RECT 7.060000 553.320000 11.820000 554.400000 ;
      RECT 0.000000 553.320000 5.260000 554.400000 ;
      RECT 0.000000 551.680000 550.160000 553.320000 ;
      RECT 547.100000 551.590000 550.160000 551.680000 ;
      RECT 547.100000 550.610000 548.960000 551.590000 ;
      RECT 547.100000 550.600000 550.160000 550.610000 ;
      RECT 506.620000 550.600000 545.300000 551.680000 ;
      RECT 461.620000 550.600000 504.820000 551.680000 ;
      RECT 416.620000 550.600000 459.820000 551.680000 ;
      RECT 371.620000 550.600000 414.820000 551.680000 ;
      RECT 326.620000 550.600000 369.820000 551.680000 ;
      RECT 281.620000 550.600000 324.820000 551.680000 ;
      RECT 236.620000 550.600000 279.820000 551.680000 ;
      RECT 191.620000 550.600000 234.820000 551.680000 ;
      RECT 146.620000 550.600000 189.820000 551.680000 ;
      RECT 101.620000 550.600000 144.820000 551.680000 ;
      RECT 56.620000 550.600000 99.820000 551.680000 ;
      RECT 11.620000 550.600000 54.820000 551.680000 ;
      RECT 4.860000 550.600000 9.655000 551.680000 ;
      RECT 0.000000 550.600000 3.060000 551.680000 ;
      RECT 0.000000 548.960000 550.160000 550.600000 ;
      RECT 544.900000 548.540000 550.160000 548.960000 ;
      RECT 544.900000 547.880000 548.960000 548.540000 ;
      RECT 508.620000 547.880000 543.100000 548.960000 ;
      RECT 463.620000 547.880000 506.820000 548.960000 ;
      RECT 418.620000 547.880000 461.820000 548.960000 ;
      RECT 373.620000 547.880000 416.820000 548.960000 ;
      RECT 328.620000 547.880000 371.820000 548.960000 ;
      RECT 283.620000 547.880000 326.820000 548.960000 ;
      RECT 238.620000 547.880000 281.820000 548.960000 ;
      RECT 193.620000 547.880000 236.820000 548.960000 ;
      RECT 148.620000 547.880000 191.820000 548.960000 ;
      RECT 103.620000 547.880000 146.820000 548.960000 ;
      RECT 58.620000 547.880000 101.820000 548.960000 ;
      RECT 13.620000 547.880000 56.820000 548.960000 ;
      RECT 7.060000 547.880000 11.820000 548.960000 ;
      RECT 0.000000 547.880000 5.260000 548.960000 ;
      RECT 0.000000 547.560000 548.960000 547.880000 ;
      RECT 0.000000 546.240000 550.160000 547.560000 ;
      RECT 547.100000 545.160000 550.160000 546.240000 ;
      RECT 506.620000 545.160000 545.300000 546.240000 ;
      RECT 461.620000 545.160000 504.820000 546.240000 ;
      RECT 416.620000 545.160000 459.820000 546.240000 ;
      RECT 371.620000 545.160000 414.820000 546.240000 ;
      RECT 326.620000 545.160000 369.820000 546.240000 ;
      RECT 281.620000 545.160000 324.820000 546.240000 ;
      RECT 236.620000 545.160000 279.820000 546.240000 ;
      RECT 191.620000 545.160000 234.820000 546.240000 ;
      RECT 146.620000 545.160000 189.820000 546.240000 ;
      RECT 101.620000 545.160000 144.820000 546.240000 ;
      RECT 56.620000 545.160000 99.820000 546.240000 ;
      RECT 11.620000 545.160000 54.820000 546.240000 ;
      RECT 4.860000 545.160000 9.655000 546.240000 ;
      RECT 0.000000 545.160000 3.060000 546.240000 ;
      RECT 0.000000 544.880000 550.160000 545.160000 ;
      RECT 0.000000 543.900000 548.960000 544.880000 ;
      RECT 0.000000 543.520000 550.160000 543.900000 ;
      RECT 544.900000 542.440000 550.160000 543.520000 ;
      RECT 508.620000 542.440000 543.100000 543.520000 ;
      RECT 463.620000 542.440000 506.820000 543.520000 ;
      RECT 418.620000 542.440000 461.820000 543.520000 ;
      RECT 373.620000 542.440000 416.820000 543.520000 ;
      RECT 328.620000 542.440000 371.820000 543.520000 ;
      RECT 283.620000 542.440000 326.820000 543.520000 ;
      RECT 238.620000 542.440000 281.820000 543.520000 ;
      RECT 193.620000 542.440000 236.820000 543.520000 ;
      RECT 148.620000 542.440000 191.820000 543.520000 ;
      RECT 103.620000 542.440000 146.820000 543.520000 ;
      RECT 58.620000 542.440000 101.820000 543.520000 ;
      RECT 13.620000 542.440000 56.820000 543.520000 ;
      RECT 7.060000 542.440000 11.820000 543.520000 ;
      RECT 0.000000 542.440000 5.260000 543.520000 ;
      RECT 0.000000 541.220000 550.160000 542.440000 ;
      RECT 0.000000 540.800000 548.960000 541.220000 ;
      RECT 547.100000 540.240000 548.960000 540.800000 ;
      RECT 547.100000 539.720000 550.160000 540.240000 ;
      RECT 506.620000 539.720000 545.300000 540.800000 ;
      RECT 461.620000 539.720000 504.820000 540.800000 ;
      RECT 416.620000 539.720000 459.820000 540.800000 ;
      RECT 371.620000 539.720000 414.820000 540.800000 ;
      RECT 326.620000 539.720000 369.820000 540.800000 ;
      RECT 281.620000 539.720000 324.820000 540.800000 ;
      RECT 236.620000 539.720000 279.820000 540.800000 ;
      RECT 191.620000 539.720000 234.820000 540.800000 ;
      RECT 146.620000 539.720000 189.820000 540.800000 ;
      RECT 101.620000 539.720000 144.820000 540.800000 ;
      RECT 56.620000 539.720000 99.820000 540.800000 ;
      RECT 11.620000 539.720000 54.820000 540.800000 ;
      RECT 4.860000 539.720000 9.655000 540.800000 ;
      RECT 0.000000 539.720000 3.060000 540.800000 ;
      RECT 0.000000 538.170000 550.160000 539.720000 ;
      RECT 0.000000 538.080000 548.960000 538.170000 ;
      RECT 544.900000 537.190000 548.960000 538.080000 ;
      RECT 544.900000 537.000000 550.160000 537.190000 ;
      RECT 508.620000 537.000000 543.100000 538.080000 ;
      RECT 463.620000 537.000000 506.820000 538.080000 ;
      RECT 418.620000 537.000000 461.820000 538.080000 ;
      RECT 373.620000 537.000000 416.820000 538.080000 ;
      RECT 328.620000 537.000000 371.820000 538.080000 ;
      RECT 283.620000 537.000000 326.820000 538.080000 ;
      RECT 238.620000 537.000000 281.820000 538.080000 ;
      RECT 193.620000 537.000000 236.820000 538.080000 ;
      RECT 148.620000 537.000000 191.820000 538.080000 ;
      RECT 103.620000 537.000000 146.820000 538.080000 ;
      RECT 58.620000 537.000000 101.820000 538.080000 ;
      RECT 13.620000 537.000000 56.820000 538.080000 ;
      RECT 7.060000 537.000000 11.820000 538.080000 ;
      RECT 0.000000 537.000000 5.260000 538.080000 ;
      RECT 0.000000 535.360000 550.160000 537.000000 ;
      RECT 547.100000 534.510000 550.160000 535.360000 ;
      RECT 547.100000 534.280000 548.960000 534.510000 ;
      RECT 506.620000 534.280000 545.300000 535.360000 ;
      RECT 461.620000 534.280000 504.820000 535.360000 ;
      RECT 416.620000 534.280000 459.820000 535.360000 ;
      RECT 371.620000 534.280000 414.820000 535.360000 ;
      RECT 326.620000 534.280000 369.820000 535.360000 ;
      RECT 281.620000 534.280000 324.820000 535.360000 ;
      RECT 236.620000 534.280000 279.820000 535.360000 ;
      RECT 191.620000 534.280000 234.820000 535.360000 ;
      RECT 146.620000 534.280000 189.820000 535.360000 ;
      RECT 101.620000 534.280000 144.820000 535.360000 ;
      RECT 56.620000 534.280000 99.820000 535.360000 ;
      RECT 11.620000 534.280000 54.820000 535.360000 ;
      RECT 4.860000 534.280000 9.655000 535.360000 ;
      RECT 0.000000 534.280000 3.060000 535.360000 ;
      RECT 0.000000 533.530000 548.960000 534.280000 ;
      RECT 0.000000 532.640000 550.160000 533.530000 ;
      RECT 544.900000 531.560000 550.160000 532.640000 ;
      RECT 508.620000 531.560000 543.100000 532.640000 ;
      RECT 463.620000 531.560000 506.820000 532.640000 ;
      RECT 418.620000 531.560000 461.820000 532.640000 ;
      RECT 373.620000 531.560000 416.820000 532.640000 ;
      RECT 328.620000 531.560000 371.820000 532.640000 ;
      RECT 283.620000 531.560000 326.820000 532.640000 ;
      RECT 238.620000 531.560000 281.820000 532.640000 ;
      RECT 193.620000 531.560000 236.820000 532.640000 ;
      RECT 148.620000 531.560000 191.820000 532.640000 ;
      RECT 103.620000 531.560000 146.820000 532.640000 ;
      RECT 58.620000 531.560000 101.820000 532.640000 ;
      RECT 13.620000 531.560000 56.820000 532.640000 ;
      RECT 7.060000 531.560000 11.820000 532.640000 ;
      RECT 0.000000 531.560000 5.260000 532.640000 ;
      RECT 0.000000 530.850000 550.160000 531.560000 ;
      RECT 0.000000 529.920000 548.960000 530.850000 ;
      RECT 547.100000 529.870000 548.960000 529.920000 ;
      RECT 547.100000 528.840000 550.160000 529.870000 ;
      RECT 506.620000 528.840000 545.300000 529.920000 ;
      RECT 461.620000 528.840000 504.820000 529.920000 ;
      RECT 416.620000 528.840000 459.820000 529.920000 ;
      RECT 371.620000 528.840000 414.820000 529.920000 ;
      RECT 326.620000 528.840000 369.820000 529.920000 ;
      RECT 281.620000 528.840000 324.820000 529.920000 ;
      RECT 236.620000 528.840000 279.820000 529.920000 ;
      RECT 191.620000 528.840000 234.820000 529.920000 ;
      RECT 146.620000 528.840000 189.820000 529.920000 ;
      RECT 101.620000 528.840000 144.820000 529.920000 ;
      RECT 56.620000 528.840000 99.820000 529.920000 ;
      RECT 11.620000 528.840000 54.820000 529.920000 ;
      RECT 4.860000 528.840000 9.655000 529.920000 ;
      RECT 0.000000 528.840000 3.060000 529.920000 ;
      RECT 0.000000 527.800000 550.160000 528.840000 ;
      RECT 0.000000 527.200000 548.960000 527.800000 ;
      RECT 544.900000 526.820000 548.960000 527.200000 ;
      RECT 544.900000 526.120000 550.160000 526.820000 ;
      RECT 508.620000 526.120000 543.100000 527.200000 ;
      RECT 463.620000 526.120000 506.820000 527.200000 ;
      RECT 418.620000 526.120000 461.820000 527.200000 ;
      RECT 373.620000 526.120000 416.820000 527.200000 ;
      RECT 328.620000 526.120000 371.820000 527.200000 ;
      RECT 283.620000 526.120000 326.820000 527.200000 ;
      RECT 238.620000 526.120000 281.820000 527.200000 ;
      RECT 193.620000 526.120000 236.820000 527.200000 ;
      RECT 148.620000 526.120000 191.820000 527.200000 ;
      RECT 103.620000 526.120000 146.820000 527.200000 ;
      RECT 58.620000 526.120000 101.820000 527.200000 ;
      RECT 13.620000 526.120000 56.820000 527.200000 ;
      RECT 7.060000 526.120000 11.820000 527.200000 ;
      RECT 0.000000 526.120000 5.260000 527.200000 ;
      RECT 0.000000 524.480000 550.160000 526.120000 ;
      RECT 547.100000 524.140000 550.160000 524.480000 ;
      RECT 547.100000 523.400000 548.960000 524.140000 ;
      RECT 506.620000 523.400000 545.300000 524.480000 ;
      RECT 461.620000 523.400000 504.820000 524.480000 ;
      RECT 416.620000 523.400000 459.820000 524.480000 ;
      RECT 371.620000 523.400000 414.820000 524.480000 ;
      RECT 326.620000 523.400000 369.820000 524.480000 ;
      RECT 281.620000 523.400000 324.820000 524.480000 ;
      RECT 236.620000 523.400000 279.820000 524.480000 ;
      RECT 191.620000 523.400000 234.820000 524.480000 ;
      RECT 146.620000 523.400000 189.820000 524.480000 ;
      RECT 101.620000 523.400000 144.820000 524.480000 ;
      RECT 56.620000 523.400000 99.820000 524.480000 ;
      RECT 11.620000 523.400000 54.820000 524.480000 ;
      RECT 4.860000 523.400000 9.655000 524.480000 ;
      RECT 0.000000 523.400000 3.060000 524.480000 ;
      RECT 0.000000 523.160000 548.960000 523.400000 ;
      RECT 0.000000 521.760000 550.160000 523.160000 ;
      RECT 544.900000 520.680000 550.160000 521.760000 ;
      RECT 508.620000 520.680000 543.100000 521.760000 ;
      RECT 463.620000 520.680000 506.820000 521.760000 ;
      RECT 418.620000 520.680000 461.820000 521.760000 ;
      RECT 373.620000 520.680000 416.820000 521.760000 ;
      RECT 328.620000 520.680000 371.820000 521.760000 ;
      RECT 283.620000 520.680000 326.820000 521.760000 ;
      RECT 238.620000 520.680000 281.820000 521.760000 ;
      RECT 193.620000 520.680000 236.820000 521.760000 ;
      RECT 148.620000 520.680000 191.820000 521.760000 ;
      RECT 103.620000 520.680000 146.820000 521.760000 ;
      RECT 58.620000 520.680000 101.820000 521.760000 ;
      RECT 13.620000 520.680000 56.820000 521.760000 ;
      RECT 7.060000 520.680000 11.820000 521.760000 ;
      RECT 0.000000 520.680000 5.260000 521.760000 ;
      RECT 0.000000 520.480000 550.160000 520.680000 ;
      RECT 0.000000 519.500000 548.960000 520.480000 ;
      RECT 0.000000 519.040000 550.160000 519.500000 ;
      RECT 547.100000 517.960000 550.160000 519.040000 ;
      RECT 506.620000 517.960000 545.300000 519.040000 ;
      RECT 461.620000 517.960000 504.820000 519.040000 ;
      RECT 416.620000 517.960000 459.820000 519.040000 ;
      RECT 371.620000 517.960000 414.820000 519.040000 ;
      RECT 326.620000 517.960000 369.820000 519.040000 ;
      RECT 281.620000 517.960000 324.820000 519.040000 ;
      RECT 236.620000 517.960000 279.820000 519.040000 ;
      RECT 191.620000 517.960000 234.820000 519.040000 ;
      RECT 146.620000 517.960000 189.820000 519.040000 ;
      RECT 101.620000 517.960000 144.820000 519.040000 ;
      RECT 56.620000 517.960000 99.820000 519.040000 ;
      RECT 11.620000 517.960000 54.820000 519.040000 ;
      RECT 4.860000 517.960000 9.655000 519.040000 ;
      RECT 0.000000 517.960000 3.060000 519.040000 ;
      RECT 0.000000 517.430000 550.160000 517.960000 ;
      RECT 0.000000 516.450000 548.960000 517.430000 ;
      RECT 0.000000 516.320000 550.160000 516.450000 ;
      RECT 544.900000 515.240000 550.160000 516.320000 ;
      RECT 508.620000 515.240000 543.100000 516.320000 ;
      RECT 463.620000 515.240000 506.820000 516.320000 ;
      RECT 418.620000 515.240000 461.820000 516.320000 ;
      RECT 373.620000 515.240000 416.820000 516.320000 ;
      RECT 328.620000 515.240000 371.820000 516.320000 ;
      RECT 283.620000 515.240000 326.820000 516.320000 ;
      RECT 238.620000 515.240000 281.820000 516.320000 ;
      RECT 193.620000 515.240000 236.820000 516.320000 ;
      RECT 148.620000 515.240000 191.820000 516.320000 ;
      RECT 103.620000 515.240000 146.820000 516.320000 ;
      RECT 58.620000 515.240000 101.820000 516.320000 ;
      RECT 13.620000 515.240000 56.820000 516.320000 ;
      RECT 7.060000 515.240000 11.820000 516.320000 ;
      RECT 0.000000 515.240000 5.260000 516.320000 ;
      RECT 0.000000 513.770000 550.160000 515.240000 ;
      RECT 0.000000 513.600000 548.960000 513.770000 ;
      RECT 547.100000 512.790000 548.960000 513.600000 ;
      RECT 547.100000 512.520000 550.160000 512.790000 ;
      RECT 506.620000 512.520000 545.300000 513.600000 ;
      RECT 461.620000 512.520000 504.820000 513.600000 ;
      RECT 416.620000 512.520000 459.820000 513.600000 ;
      RECT 371.620000 512.520000 414.820000 513.600000 ;
      RECT 326.620000 512.520000 369.820000 513.600000 ;
      RECT 281.620000 512.520000 324.820000 513.600000 ;
      RECT 236.620000 512.520000 279.820000 513.600000 ;
      RECT 191.620000 512.520000 234.820000 513.600000 ;
      RECT 146.620000 512.520000 189.820000 513.600000 ;
      RECT 101.620000 512.520000 144.820000 513.600000 ;
      RECT 56.620000 512.520000 99.820000 513.600000 ;
      RECT 11.620000 512.520000 54.820000 513.600000 ;
      RECT 4.860000 512.520000 9.655000 513.600000 ;
      RECT 0.000000 512.520000 3.060000 513.600000 ;
      RECT 0.000000 510.880000 550.160000 512.520000 ;
      RECT 544.900000 510.110000 550.160000 510.880000 ;
      RECT 544.900000 509.800000 548.960000 510.110000 ;
      RECT 508.620000 509.800000 543.100000 510.880000 ;
      RECT 463.620000 509.800000 506.820000 510.880000 ;
      RECT 418.620000 509.800000 461.820000 510.880000 ;
      RECT 373.620000 509.800000 416.820000 510.880000 ;
      RECT 328.620000 509.800000 371.820000 510.880000 ;
      RECT 283.620000 509.800000 326.820000 510.880000 ;
      RECT 238.620000 509.800000 281.820000 510.880000 ;
      RECT 193.620000 509.800000 236.820000 510.880000 ;
      RECT 148.620000 509.800000 191.820000 510.880000 ;
      RECT 103.620000 509.800000 146.820000 510.880000 ;
      RECT 58.620000 509.800000 101.820000 510.880000 ;
      RECT 13.620000 509.800000 56.820000 510.880000 ;
      RECT 7.060000 509.800000 11.820000 510.880000 ;
      RECT 0.000000 509.800000 5.260000 510.880000 ;
      RECT 0.000000 509.130000 548.960000 509.800000 ;
      RECT 0.000000 508.160000 550.160000 509.130000 ;
      RECT 547.100000 507.080000 550.160000 508.160000 ;
      RECT 506.620000 507.080000 545.300000 508.160000 ;
      RECT 461.620000 507.080000 504.820000 508.160000 ;
      RECT 416.620000 507.080000 459.820000 508.160000 ;
      RECT 371.620000 507.080000 414.820000 508.160000 ;
      RECT 326.620000 507.080000 369.820000 508.160000 ;
      RECT 281.620000 507.080000 324.820000 508.160000 ;
      RECT 236.620000 507.080000 279.820000 508.160000 ;
      RECT 191.620000 507.080000 234.820000 508.160000 ;
      RECT 146.620000 507.080000 189.820000 508.160000 ;
      RECT 101.620000 507.080000 144.820000 508.160000 ;
      RECT 56.620000 507.080000 99.820000 508.160000 ;
      RECT 11.620000 507.080000 54.820000 508.160000 ;
      RECT 4.860000 507.080000 9.655000 508.160000 ;
      RECT 0.000000 507.080000 3.060000 508.160000 ;
      RECT 0.000000 507.060000 550.160000 507.080000 ;
      RECT 0.000000 506.080000 548.960000 507.060000 ;
      RECT 0.000000 505.440000 550.160000 506.080000 ;
      RECT 544.900000 504.360000 550.160000 505.440000 ;
      RECT 508.620000 504.360000 543.100000 505.440000 ;
      RECT 463.620000 504.360000 506.820000 505.440000 ;
      RECT 418.620000 504.360000 461.820000 505.440000 ;
      RECT 373.620000 504.360000 416.820000 505.440000 ;
      RECT 328.620000 504.360000 371.820000 505.440000 ;
      RECT 283.620000 504.360000 326.820000 505.440000 ;
      RECT 238.620000 504.360000 281.820000 505.440000 ;
      RECT 193.620000 504.360000 236.820000 505.440000 ;
      RECT 148.620000 504.360000 191.820000 505.440000 ;
      RECT 103.620000 504.360000 146.820000 505.440000 ;
      RECT 58.620000 504.360000 101.820000 505.440000 ;
      RECT 13.620000 504.360000 56.820000 505.440000 ;
      RECT 7.060000 504.360000 11.820000 505.440000 ;
      RECT 0.000000 504.360000 5.260000 505.440000 ;
      RECT 0.000000 503.400000 550.160000 504.360000 ;
      RECT 0.000000 502.720000 548.960000 503.400000 ;
      RECT 547.100000 502.420000 548.960000 502.720000 ;
      RECT 547.100000 501.640000 550.160000 502.420000 ;
      RECT 506.620000 501.640000 545.300000 502.720000 ;
      RECT 461.620000 501.640000 504.820000 502.720000 ;
      RECT 416.620000 501.640000 459.820000 502.720000 ;
      RECT 371.620000 501.640000 414.820000 502.720000 ;
      RECT 326.620000 501.640000 369.820000 502.720000 ;
      RECT 281.620000 501.640000 324.820000 502.720000 ;
      RECT 236.620000 501.640000 279.820000 502.720000 ;
      RECT 191.620000 501.640000 234.820000 502.720000 ;
      RECT 146.620000 501.640000 189.820000 502.720000 ;
      RECT 101.620000 501.640000 144.820000 502.720000 ;
      RECT 56.620000 501.640000 99.820000 502.720000 ;
      RECT 11.620000 501.640000 54.820000 502.720000 ;
      RECT 4.860000 501.640000 9.655000 502.720000 ;
      RECT 0.000000 501.640000 3.060000 502.720000 ;
      RECT 0.000000 500.000000 550.160000 501.640000 ;
      RECT 544.900000 499.740000 550.160000 500.000000 ;
      RECT 544.900000 498.920000 548.960000 499.740000 ;
      RECT 508.620000 498.920000 543.100000 500.000000 ;
      RECT 463.620000 498.920000 506.820000 500.000000 ;
      RECT 418.620000 498.920000 461.820000 500.000000 ;
      RECT 373.620000 498.920000 416.820000 500.000000 ;
      RECT 328.620000 498.920000 371.820000 500.000000 ;
      RECT 283.620000 498.920000 326.820000 500.000000 ;
      RECT 238.620000 498.920000 281.820000 500.000000 ;
      RECT 193.620000 498.920000 236.820000 500.000000 ;
      RECT 148.620000 498.920000 191.820000 500.000000 ;
      RECT 103.620000 498.920000 146.820000 500.000000 ;
      RECT 58.620000 498.920000 101.820000 500.000000 ;
      RECT 13.620000 498.920000 56.820000 500.000000 ;
      RECT 7.060000 498.920000 11.820000 500.000000 ;
      RECT 0.000000 498.920000 5.260000 500.000000 ;
      RECT 0.000000 498.760000 548.960000 498.920000 ;
      RECT 0.000000 497.280000 550.160000 498.760000 ;
      RECT 547.100000 496.690000 550.160000 497.280000 ;
      RECT 547.100000 496.200000 548.960000 496.690000 ;
      RECT 506.620000 496.200000 545.300000 497.280000 ;
      RECT 461.620000 496.200000 504.820000 497.280000 ;
      RECT 416.620000 496.200000 459.820000 497.280000 ;
      RECT 371.620000 496.200000 414.820000 497.280000 ;
      RECT 326.620000 496.200000 369.820000 497.280000 ;
      RECT 281.620000 496.200000 324.820000 497.280000 ;
      RECT 236.620000 496.200000 279.820000 497.280000 ;
      RECT 191.620000 496.200000 234.820000 497.280000 ;
      RECT 146.620000 496.200000 189.820000 497.280000 ;
      RECT 101.620000 496.200000 144.820000 497.280000 ;
      RECT 56.620000 496.200000 99.820000 497.280000 ;
      RECT 11.620000 496.200000 54.820000 497.280000 ;
      RECT 4.860000 496.200000 9.655000 497.280000 ;
      RECT 0.000000 496.200000 3.060000 497.280000 ;
      RECT 0.000000 495.710000 548.960000 496.200000 ;
      RECT 0.000000 494.560000 550.160000 495.710000 ;
      RECT 544.900000 493.480000 550.160000 494.560000 ;
      RECT 508.620000 493.480000 543.100000 494.560000 ;
      RECT 463.620000 493.480000 506.820000 494.560000 ;
      RECT 418.620000 493.480000 461.820000 494.560000 ;
      RECT 373.620000 493.480000 416.820000 494.560000 ;
      RECT 328.620000 493.480000 371.820000 494.560000 ;
      RECT 283.620000 493.480000 326.820000 494.560000 ;
      RECT 238.620000 493.480000 281.820000 494.560000 ;
      RECT 193.620000 493.480000 236.820000 494.560000 ;
      RECT 148.620000 493.480000 191.820000 494.560000 ;
      RECT 103.620000 493.480000 146.820000 494.560000 ;
      RECT 58.620000 493.480000 101.820000 494.560000 ;
      RECT 13.620000 493.480000 56.820000 494.560000 ;
      RECT 7.060000 493.480000 11.820000 494.560000 ;
      RECT 0.000000 493.480000 5.260000 494.560000 ;
      RECT 0.000000 493.030000 550.160000 493.480000 ;
      RECT 0.000000 492.050000 548.960000 493.030000 ;
      RECT 0.000000 491.840000 550.160000 492.050000 ;
      RECT 547.100000 490.760000 550.160000 491.840000 ;
      RECT 506.620000 490.760000 545.300000 491.840000 ;
      RECT 461.620000 490.760000 504.820000 491.840000 ;
      RECT 416.620000 490.760000 459.820000 491.840000 ;
      RECT 371.620000 490.760000 414.820000 491.840000 ;
      RECT 326.620000 490.760000 369.820000 491.840000 ;
      RECT 281.620000 490.760000 324.820000 491.840000 ;
      RECT 236.620000 490.760000 279.820000 491.840000 ;
      RECT 191.620000 490.760000 234.820000 491.840000 ;
      RECT 146.620000 490.760000 189.820000 491.840000 ;
      RECT 101.620000 490.760000 144.820000 491.840000 ;
      RECT 56.620000 490.760000 99.820000 491.840000 ;
      RECT 11.620000 490.760000 54.820000 491.840000 ;
      RECT 4.860000 490.760000 9.655000 491.840000 ;
      RECT 0.000000 490.760000 3.060000 491.840000 ;
      RECT 0.000000 489.980000 550.160000 490.760000 ;
      RECT 0.000000 489.120000 548.960000 489.980000 ;
      RECT 544.900000 489.000000 548.960000 489.120000 ;
      RECT 544.900000 488.040000 550.160000 489.000000 ;
      RECT 508.620000 488.040000 543.100000 489.120000 ;
      RECT 463.620000 488.040000 506.820000 489.120000 ;
      RECT 418.620000 488.040000 461.820000 489.120000 ;
      RECT 373.620000 488.040000 416.820000 489.120000 ;
      RECT 328.620000 488.040000 371.820000 489.120000 ;
      RECT 283.620000 488.040000 326.820000 489.120000 ;
      RECT 238.620000 488.040000 281.820000 489.120000 ;
      RECT 193.620000 488.040000 236.820000 489.120000 ;
      RECT 148.620000 488.040000 191.820000 489.120000 ;
      RECT 103.620000 488.040000 146.820000 489.120000 ;
      RECT 58.620000 488.040000 101.820000 489.120000 ;
      RECT 13.620000 488.040000 56.820000 489.120000 ;
      RECT 7.060000 488.040000 11.820000 489.120000 ;
      RECT 0.000000 488.040000 5.260000 489.120000 ;
      RECT 0.000000 486.400000 550.160000 488.040000 ;
      RECT 547.100000 486.320000 550.160000 486.400000 ;
      RECT 547.100000 485.340000 548.960000 486.320000 ;
      RECT 547.100000 485.320000 550.160000 485.340000 ;
      RECT 506.620000 485.320000 545.300000 486.400000 ;
      RECT 461.620000 485.320000 504.820000 486.400000 ;
      RECT 416.620000 485.320000 459.820000 486.400000 ;
      RECT 371.620000 485.320000 414.820000 486.400000 ;
      RECT 326.620000 485.320000 369.820000 486.400000 ;
      RECT 281.620000 485.320000 324.820000 486.400000 ;
      RECT 236.620000 485.320000 279.820000 486.400000 ;
      RECT 191.620000 485.320000 234.820000 486.400000 ;
      RECT 146.620000 485.320000 189.820000 486.400000 ;
      RECT 101.620000 485.320000 144.820000 486.400000 ;
      RECT 56.620000 485.320000 99.820000 486.400000 ;
      RECT 11.620000 485.320000 54.820000 486.400000 ;
      RECT 4.860000 485.320000 9.655000 486.400000 ;
      RECT 0.000000 485.320000 3.060000 486.400000 ;
      RECT 0.000000 483.680000 550.160000 485.320000 ;
      RECT 544.900000 482.660000 550.160000 483.680000 ;
      RECT 544.900000 482.600000 548.960000 482.660000 ;
      RECT 508.620000 482.600000 543.100000 483.680000 ;
      RECT 463.620000 482.600000 506.820000 483.680000 ;
      RECT 418.620000 482.600000 461.820000 483.680000 ;
      RECT 373.620000 482.600000 416.820000 483.680000 ;
      RECT 328.620000 482.600000 371.820000 483.680000 ;
      RECT 283.620000 482.600000 326.820000 483.680000 ;
      RECT 238.620000 482.600000 281.820000 483.680000 ;
      RECT 193.620000 482.600000 236.820000 483.680000 ;
      RECT 148.620000 482.600000 191.820000 483.680000 ;
      RECT 103.620000 482.600000 146.820000 483.680000 ;
      RECT 58.620000 482.600000 101.820000 483.680000 ;
      RECT 13.620000 482.600000 56.820000 483.680000 ;
      RECT 7.060000 482.600000 11.820000 483.680000 ;
      RECT 0.000000 482.600000 5.260000 483.680000 ;
      RECT 0.000000 481.680000 548.960000 482.600000 ;
      RECT 0.000000 480.960000 550.160000 481.680000 ;
      RECT 547.100000 479.880000 550.160000 480.960000 ;
      RECT 506.620000 479.880000 545.300000 480.960000 ;
      RECT 461.620000 479.880000 504.820000 480.960000 ;
      RECT 416.620000 479.880000 459.820000 480.960000 ;
      RECT 371.620000 479.880000 414.820000 480.960000 ;
      RECT 326.620000 479.880000 369.820000 480.960000 ;
      RECT 281.620000 479.880000 324.820000 480.960000 ;
      RECT 236.620000 479.880000 279.820000 480.960000 ;
      RECT 191.620000 479.880000 234.820000 480.960000 ;
      RECT 146.620000 479.880000 189.820000 480.960000 ;
      RECT 101.620000 479.880000 144.820000 480.960000 ;
      RECT 56.620000 479.880000 99.820000 480.960000 ;
      RECT 11.620000 479.880000 54.820000 480.960000 ;
      RECT 4.860000 479.880000 9.655000 480.960000 ;
      RECT 0.000000 479.880000 3.060000 480.960000 ;
      RECT 0.000000 479.610000 550.160000 479.880000 ;
      RECT 0.000000 478.630000 548.960000 479.610000 ;
      RECT 0.000000 478.240000 550.160000 478.630000 ;
      RECT 544.900000 477.160000 550.160000 478.240000 ;
      RECT 508.620000 477.160000 543.100000 478.240000 ;
      RECT 463.620000 477.160000 506.820000 478.240000 ;
      RECT 418.620000 477.160000 461.820000 478.240000 ;
      RECT 373.620000 477.160000 416.820000 478.240000 ;
      RECT 328.620000 477.160000 371.820000 478.240000 ;
      RECT 283.620000 477.160000 326.820000 478.240000 ;
      RECT 238.620000 477.160000 281.820000 478.240000 ;
      RECT 193.620000 477.160000 236.820000 478.240000 ;
      RECT 148.620000 477.160000 191.820000 478.240000 ;
      RECT 103.620000 477.160000 146.820000 478.240000 ;
      RECT 58.620000 477.160000 101.820000 478.240000 ;
      RECT 13.620000 477.160000 56.820000 478.240000 ;
      RECT 7.060000 477.160000 11.820000 478.240000 ;
      RECT 0.000000 477.160000 5.260000 478.240000 ;
      RECT 0.000000 475.950000 550.160000 477.160000 ;
      RECT 0.000000 475.520000 548.960000 475.950000 ;
      RECT 547.100000 474.970000 548.960000 475.520000 ;
      RECT 547.100000 474.440000 550.160000 474.970000 ;
      RECT 506.620000 474.440000 545.300000 475.520000 ;
      RECT 461.620000 474.440000 504.820000 475.520000 ;
      RECT 416.620000 474.440000 459.820000 475.520000 ;
      RECT 371.620000 474.440000 414.820000 475.520000 ;
      RECT 326.620000 474.440000 369.820000 475.520000 ;
      RECT 281.620000 474.440000 324.820000 475.520000 ;
      RECT 236.620000 474.440000 279.820000 475.520000 ;
      RECT 191.620000 474.440000 234.820000 475.520000 ;
      RECT 146.620000 474.440000 189.820000 475.520000 ;
      RECT 101.620000 474.440000 144.820000 475.520000 ;
      RECT 56.620000 474.440000 99.820000 475.520000 ;
      RECT 11.620000 474.440000 54.820000 475.520000 ;
      RECT 4.860000 474.440000 9.655000 475.520000 ;
      RECT 0.000000 474.440000 3.060000 475.520000 ;
      RECT 0.000000 472.800000 550.160000 474.440000 ;
      RECT 544.900000 472.290000 550.160000 472.800000 ;
      RECT 544.900000 471.720000 548.960000 472.290000 ;
      RECT 508.620000 471.720000 543.100000 472.800000 ;
      RECT 463.620000 471.720000 506.820000 472.800000 ;
      RECT 418.620000 471.720000 461.820000 472.800000 ;
      RECT 373.620000 471.720000 416.820000 472.800000 ;
      RECT 328.620000 471.720000 371.820000 472.800000 ;
      RECT 283.620000 471.720000 326.820000 472.800000 ;
      RECT 238.620000 471.720000 281.820000 472.800000 ;
      RECT 193.620000 471.720000 236.820000 472.800000 ;
      RECT 148.620000 471.720000 191.820000 472.800000 ;
      RECT 103.620000 471.720000 146.820000 472.800000 ;
      RECT 58.620000 471.720000 101.820000 472.800000 ;
      RECT 13.620000 471.720000 56.820000 472.800000 ;
      RECT 7.060000 471.720000 11.820000 472.800000 ;
      RECT 0.000000 471.720000 5.260000 472.800000 ;
      RECT 0.000000 471.310000 548.960000 471.720000 ;
      RECT 0.000000 470.080000 550.160000 471.310000 ;
      RECT 547.100000 469.240000 550.160000 470.080000 ;
      RECT 547.100000 469.000000 548.960000 469.240000 ;
      RECT 506.620000 469.000000 545.300000 470.080000 ;
      RECT 461.620000 469.000000 504.820000 470.080000 ;
      RECT 416.620000 469.000000 459.820000 470.080000 ;
      RECT 371.620000 469.000000 414.820000 470.080000 ;
      RECT 326.620000 469.000000 369.820000 470.080000 ;
      RECT 281.620000 469.000000 324.820000 470.080000 ;
      RECT 236.620000 469.000000 279.820000 470.080000 ;
      RECT 191.620000 469.000000 234.820000 470.080000 ;
      RECT 146.620000 469.000000 189.820000 470.080000 ;
      RECT 101.620000 469.000000 144.820000 470.080000 ;
      RECT 56.620000 469.000000 99.820000 470.080000 ;
      RECT 11.620000 469.000000 54.820000 470.080000 ;
      RECT 4.860000 469.000000 9.655000 470.080000 ;
      RECT 0.000000 469.000000 3.060000 470.080000 ;
      RECT 0.000000 468.260000 548.960000 469.000000 ;
      RECT 0.000000 467.360000 550.160000 468.260000 ;
      RECT 544.900000 466.280000 550.160000 467.360000 ;
      RECT 508.620000 466.280000 543.100000 467.360000 ;
      RECT 463.620000 466.280000 506.820000 467.360000 ;
      RECT 418.620000 466.280000 461.820000 467.360000 ;
      RECT 373.620000 466.280000 416.820000 467.360000 ;
      RECT 328.620000 466.280000 371.820000 467.360000 ;
      RECT 283.620000 466.280000 326.820000 467.360000 ;
      RECT 238.620000 466.280000 281.820000 467.360000 ;
      RECT 193.620000 466.280000 236.820000 467.360000 ;
      RECT 148.620000 466.280000 191.820000 467.360000 ;
      RECT 103.620000 466.280000 146.820000 467.360000 ;
      RECT 58.620000 466.280000 101.820000 467.360000 ;
      RECT 13.620000 466.280000 56.820000 467.360000 ;
      RECT 7.060000 466.280000 11.820000 467.360000 ;
      RECT 0.000000 466.280000 5.260000 467.360000 ;
      RECT 0.000000 465.580000 550.160000 466.280000 ;
      RECT 0.000000 464.640000 548.960000 465.580000 ;
      RECT 547.100000 464.600000 548.960000 464.640000 ;
      RECT 547.100000 463.560000 550.160000 464.600000 ;
      RECT 506.620000 463.560000 545.300000 464.640000 ;
      RECT 461.620000 463.560000 504.820000 464.640000 ;
      RECT 416.620000 463.560000 459.820000 464.640000 ;
      RECT 371.620000 463.560000 414.820000 464.640000 ;
      RECT 326.620000 463.560000 369.820000 464.640000 ;
      RECT 281.620000 463.560000 324.820000 464.640000 ;
      RECT 236.620000 463.560000 279.820000 464.640000 ;
      RECT 191.620000 463.560000 234.820000 464.640000 ;
      RECT 146.620000 463.560000 189.820000 464.640000 ;
      RECT 101.620000 463.560000 144.820000 464.640000 ;
      RECT 56.620000 463.560000 99.820000 464.640000 ;
      RECT 11.620000 463.560000 54.820000 464.640000 ;
      RECT 4.860000 463.560000 9.655000 464.640000 ;
      RECT 0.000000 463.560000 3.060000 464.640000 ;
      RECT 0.000000 461.920000 550.160000 463.560000 ;
      RECT 544.900000 460.940000 548.960000 461.920000 ;
      RECT 544.900000 460.840000 550.160000 460.940000 ;
      RECT 508.620000 460.840000 543.100000 461.920000 ;
      RECT 463.620000 460.840000 506.820000 461.920000 ;
      RECT 418.620000 460.840000 461.820000 461.920000 ;
      RECT 373.620000 460.840000 416.820000 461.920000 ;
      RECT 328.620000 460.840000 371.820000 461.920000 ;
      RECT 283.620000 460.840000 326.820000 461.920000 ;
      RECT 238.620000 460.840000 281.820000 461.920000 ;
      RECT 193.620000 460.840000 236.820000 461.920000 ;
      RECT 148.620000 460.840000 191.820000 461.920000 ;
      RECT 103.620000 460.840000 146.820000 461.920000 ;
      RECT 58.620000 460.840000 101.820000 461.920000 ;
      RECT 13.620000 460.840000 56.820000 461.920000 ;
      RECT 7.060000 460.840000 11.820000 461.920000 ;
      RECT 0.000000 460.840000 5.260000 461.920000 ;
      RECT 0.000000 459.200000 550.160000 460.840000 ;
      RECT 547.100000 458.870000 550.160000 459.200000 ;
      RECT 547.100000 458.120000 548.960000 458.870000 ;
      RECT 506.620000 458.120000 545.300000 459.200000 ;
      RECT 461.620000 458.120000 504.820000 459.200000 ;
      RECT 416.620000 458.120000 459.820000 459.200000 ;
      RECT 371.620000 458.120000 414.820000 459.200000 ;
      RECT 326.620000 458.120000 369.820000 459.200000 ;
      RECT 281.620000 458.120000 324.820000 459.200000 ;
      RECT 236.620000 458.120000 279.820000 459.200000 ;
      RECT 191.620000 458.120000 234.820000 459.200000 ;
      RECT 146.620000 458.120000 189.820000 459.200000 ;
      RECT 101.620000 458.120000 144.820000 459.200000 ;
      RECT 56.620000 458.120000 99.820000 459.200000 ;
      RECT 11.620000 458.120000 54.820000 459.200000 ;
      RECT 4.860000 458.120000 9.655000 459.200000 ;
      RECT 0.000000 458.120000 3.060000 459.200000 ;
      RECT 0.000000 457.890000 548.960000 458.120000 ;
      RECT 0.000000 456.480000 550.160000 457.890000 ;
      RECT 544.900000 455.400000 550.160000 456.480000 ;
      RECT 508.620000 455.400000 543.100000 456.480000 ;
      RECT 463.620000 455.400000 506.820000 456.480000 ;
      RECT 418.620000 455.400000 461.820000 456.480000 ;
      RECT 373.620000 455.400000 416.820000 456.480000 ;
      RECT 328.620000 455.400000 371.820000 456.480000 ;
      RECT 283.620000 455.400000 326.820000 456.480000 ;
      RECT 238.620000 455.400000 281.820000 456.480000 ;
      RECT 193.620000 455.400000 236.820000 456.480000 ;
      RECT 148.620000 455.400000 191.820000 456.480000 ;
      RECT 103.620000 455.400000 146.820000 456.480000 ;
      RECT 58.620000 455.400000 101.820000 456.480000 ;
      RECT 13.620000 455.400000 56.820000 456.480000 ;
      RECT 7.060000 455.400000 11.820000 456.480000 ;
      RECT 0.000000 455.400000 5.260000 456.480000 ;
      RECT 0.000000 455.210000 550.160000 455.400000 ;
      RECT 0.000000 454.230000 548.960000 455.210000 ;
      RECT 0.000000 453.760000 550.160000 454.230000 ;
      RECT 547.100000 452.680000 550.160000 453.760000 ;
      RECT 506.620000 452.680000 545.300000 453.760000 ;
      RECT 461.620000 452.680000 504.820000 453.760000 ;
      RECT 416.620000 452.680000 459.820000 453.760000 ;
      RECT 371.620000 452.680000 414.820000 453.760000 ;
      RECT 326.620000 452.680000 369.820000 453.760000 ;
      RECT 281.620000 452.680000 324.820000 453.760000 ;
      RECT 236.620000 452.680000 279.820000 453.760000 ;
      RECT 191.620000 452.680000 234.820000 453.760000 ;
      RECT 146.620000 452.680000 189.820000 453.760000 ;
      RECT 101.620000 452.680000 144.820000 453.760000 ;
      RECT 56.620000 452.680000 99.820000 453.760000 ;
      RECT 11.620000 452.680000 54.820000 453.760000 ;
      RECT 4.860000 452.680000 9.655000 453.760000 ;
      RECT 0.000000 452.680000 3.060000 453.760000 ;
      RECT 0.000000 451.550000 550.160000 452.680000 ;
      RECT 0.000000 451.040000 548.960000 451.550000 ;
      RECT 544.900000 450.570000 548.960000 451.040000 ;
      RECT 544.900000 449.960000 550.160000 450.570000 ;
      RECT 508.620000 449.960000 543.100000 451.040000 ;
      RECT 463.620000 449.960000 506.820000 451.040000 ;
      RECT 418.620000 449.960000 461.820000 451.040000 ;
      RECT 373.620000 449.960000 416.820000 451.040000 ;
      RECT 328.620000 449.960000 371.820000 451.040000 ;
      RECT 283.620000 449.960000 326.820000 451.040000 ;
      RECT 238.620000 449.960000 281.820000 451.040000 ;
      RECT 193.620000 449.960000 236.820000 451.040000 ;
      RECT 148.620000 449.960000 191.820000 451.040000 ;
      RECT 103.620000 449.960000 146.820000 451.040000 ;
      RECT 58.620000 449.960000 101.820000 451.040000 ;
      RECT 13.620000 449.960000 56.820000 451.040000 ;
      RECT 7.060000 449.960000 11.820000 451.040000 ;
      RECT 0.000000 449.960000 5.260000 451.040000 ;
      RECT 0.000000 448.500000 550.160000 449.960000 ;
      RECT 0.000000 448.320000 548.960000 448.500000 ;
      RECT 547.100000 447.520000 548.960000 448.320000 ;
      RECT 547.100000 447.240000 550.160000 447.520000 ;
      RECT 506.620000 447.240000 545.300000 448.320000 ;
      RECT 461.620000 447.240000 504.820000 448.320000 ;
      RECT 416.620000 447.240000 459.820000 448.320000 ;
      RECT 371.620000 447.240000 414.820000 448.320000 ;
      RECT 326.620000 447.240000 369.820000 448.320000 ;
      RECT 281.620000 447.240000 324.820000 448.320000 ;
      RECT 236.620000 447.240000 279.820000 448.320000 ;
      RECT 191.620000 447.240000 234.820000 448.320000 ;
      RECT 146.620000 447.240000 189.820000 448.320000 ;
      RECT 101.620000 447.240000 144.820000 448.320000 ;
      RECT 56.620000 447.240000 99.820000 448.320000 ;
      RECT 11.620000 447.240000 54.820000 448.320000 ;
      RECT 4.860000 447.240000 9.655000 448.320000 ;
      RECT 0.000000 447.240000 3.060000 448.320000 ;
      RECT 0.000000 445.600000 550.160000 447.240000 ;
      RECT 544.900000 444.840000 550.160000 445.600000 ;
      RECT 544.900000 444.520000 548.960000 444.840000 ;
      RECT 508.620000 444.520000 543.100000 445.600000 ;
      RECT 463.620000 444.520000 506.820000 445.600000 ;
      RECT 418.620000 444.520000 461.820000 445.600000 ;
      RECT 373.620000 444.520000 416.820000 445.600000 ;
      RECT 328.620000 444.520000 371.820000 445.600000 ;
      RECT 283.620000 444.520000 326.820000 445.600000 ;
      RECT 238.620000 444.520000 281.820000 445.600000 ;
      RECT 193.620000 444.520000 236.820000 445.600000 ;
      RECT 148.620000 444.520000 191.820000 445.600000 ;
      RECT 103.620000 444.520000 146.820000 445.600000 ;
      RECT 58.620000 444.520000 101.820000 445.600000 ;
      RECT 13.620000 444.520000 56.820000 445.600000 ;
      RECT 7.060000 444.520000 11.820000 445.600000 ;
      RECT 0.000000 444.520000 5.260000 445.600000 ;
      RECT 0.000000 443.860000 548.960000 444.520000 ;
      RECT 0.000000 442.880000 550.160000 443.860000 ;
      RECT 547.100000 441.800000 550.160000 442.880000 ;
      RECT 506.620000 441.800000 545.300000 442.880000 ;
      RECT 461.620000 441.800000 504.820000 442.880000 ;
      RECT 416.620000 441.800000 459.820000 442.880000 ;
      RECT 371.620000 441.800000 414.820000 442.880000 ;
      RECT 326.620000 441.800000 369.820000 442.880000 ;
      RECT 281.620000 441.800000 324.820000 442.880000 ;
      RECT 236.620000 441.800000 279.820000 442.880000 ;
      RECT 191.620000 441.800000 234.820000 442.880000 ;
      RECT 146.620000 441.800000 189.820000 442.880000 ;
      RECT 101.620000 441.800000 144.820000 442.880000 ;
      RECT 56.620000 441.800000 99.820000 442.880000 ;
      RECT 11.620000 441.800000 54.820000 442.880000 ;
      RECT 4.860000 441.800000 9.655000 442.880000 ;
      RECT 0.000000 441.800000 3.060000 442.880000 ;
      RECT 0.000000 441.180000 550.160000 441.800000 ;
      RECT 0.000000 440.200000 548.960000 441.180000 ;
      RECT 0.000000 440.160000 550.160000 440.200000 ;
      RECT 544.900000 439.080000 550.160000 440.160000 ;
      RECT 508.620000 439.080000 543.100000 440.160000 ;
      RECT 463.620000 439.080000 506.820000 440.160000 ;
      RECT 418.620000 439.080000 461.820000 440.160000 ;
      RECT 373.620000 439.080000 416.820000 440.160000 ;
      RECT 328.620000 439.080000 371.820000 440.160000 ;
      RECT 283.620000 439.080000 326.820000 440.160000 ;
      RECT 238.620000 439.080000 281.820000 440.160000 ;
      RECT 193.620000 439.080000 236.820000 440.160000 ;
      RECT 148.620000 439.080000 191.820000 440.160000 ;
      RECT 103.620000 439.080000 146.820000 440.160000 ;
      RECT 58.620000 439.080000 101.820000 440.160000 ;
      RECT 13.620000 439.080000 56.820000 440.160000 ;
      RECT 7.060000 439.080000 11.820000 440.160000 ;
      RECT 0.000000 439.080000 5.260000 440.160000 ;
      RECT 0.000000 438.130000 550.160000 439.080000 ;
      RECT 0.000000 437.440000 548.960000 438.130000 ;
      RECT 547.100000 437.150000 548.960000 437.440000 ;
      RECT 547.100000 436.360000 550.160000 437.150000 ;
      RECT 506.620000 436.360000 545.300000 437.440000 ;
      RECT 461.620000 436.360000 504.820000 437.440000 ;
      RECT 416.620000 436.360000 459.820000 437.440000 ;
      RECT 371.620000 436.360000 414.820000 437.440000 ;
      RECT 326.620000 436.360000 369.820000 437.440000 ;
      RECT 281.620000 436.360000 324.820000 437.440000 ;
      RECT 236.620000 436.360000 279.820000 437.440000 ;
      RECT 191.620000 436.360000 234.820000 437.440000 ;
      RECT 146.620000 436.360000 189.820000 437.440000 ;
      RECT 101.620000 436.360000 144.820000 437.440000 ;
      RECT 56.620000 436.360000 99.820000 437.440000 ;
      RECT 11.620000 436.360000 54.820000 437.440000 ;
      RECT 4.860000 436.360000 9.655000 437.440000 ;
      RECT 0.000000 436.360000 3.060000 437.440000 ;
      RECT 0.000000 434.720000 550.160000 436.360000 ;
      RECT 544.900000 434.470000 550.160000 434.720000 ;
      RECT 544.900000 433.640000 548.960000 434.470000 ;
      RECT 508.620000 433.640000 543.100000 434.720000 ;
      RECT 463.620000 433.640000 506.820000 434.720000 ;
      RECT 418.620000 433.640000 461.820000 434.720000 ;
      RECT 373.620000 433.640000 416.820000 434.720000 ;
      RECT 328.620000 433.640000 371.820000 434.720000 ;
      RECT 283.620000 433.640000 326.820000 434.720000 ;
      RECT 238.620000 433.640000 281.820000 434.720000 ;
      RECT 193.620000 433.640000 236.820000 434.720000 ;
      RECT 148.620000 433.640000 191.820000 434.720000 ;
      RECT 103.620000 433.640000 146.820000 434.720000 ;
      RECT 58.620000 433.640000 101.820000 434.720000 ;
      RECT 13.620000 433.640000 56.820000 434.720000 ;
      RECT 7.060000 433.640000 11.820000 434.720000 ;
      RECT 0.000000 433.640000 5.260000 434.720000 ;
      RECT 0.000000 433.490000 548.960000 433.640000 ;
      RECT 0.000000 432.000000 550.160000 433.490000 ;
      RECT 547.100000 430.920000 550.160000 432.000000 ;
      RECT 506.620000 430.920000 545.300000 432.000000 ;
      RECT 461.620000 430.920000 504.820000 432.000000 ;
      RECT 416.620000 430.920000 459.820000 432.000000 ;
      RECT 371.620000 430.920000 414.820000 432.000000 ;
      RECT 326.620000 430.920000 369.820000 432.000000 ;
      RECT 281.620000 430.920000 324.820000 432.000000 ;
      RECT 236.620000 430.920000 279.820000 432.000000 ;
      RECT 191.620000 430.920000 234.820000 432.000000 ;
      RECT 146.620000 430.920000 189.820000 432.000000 ;
      RECT 101.620000 430.920000 144.820000 432.000000 ;
      RECT 56.620000 430.920000 99.820000 432.000000 ;
      RECT 11.620000 430.920000 54.820000 432.000000 ;
      RECT 4.860000 430.920000 9.655000 432.000000 ;
      RECT 0.000000 430.920000 3.060000 432.000000 ;
      RECT 0.000000 430.810000 550.160000 430.920000 ;
      RECT 0.000000 429.830000 548.960000 430.810000 ;
      RECT 0.000000 429.280000 550.160000 429.830000 ;
      RECT 544.900000 428.200000 550.160000 429.280000 ;
      RECT 508.620000 428.200000 543.100000 429.280000 ;
      RECT 463.620000 428.200000 506.820000 429.280000 ;
      RECT 418.620000 428.200000 461.820000 429.280000 ;
      RECT 373.620000 428.200000 416.820000 429.280000 ;
      RECT 328.620000 428.200000 371.820000 429.280000 ;
      RECT 283.620000 428.200000 326.820000 429.280000 ;
      RECT 238.620000 428.200000 281.820000 429.280000 ;
      RECT 193.620000 428.200000 236.820000 429.280000 ;
      RECT 148.620000 428.200000 191.820000 429.280000 ;
      RECT 103.620000 428.200000 146.820000 429.280000 ;
      RECT 58.620000 428.200000 101.820000 429.280000 ;
      RECT 13.620000 428.200000 56.820000 429.280000 ;
      RECT 7.060000 428.200000 11.820000 429.280000 ;
      RECT 0.000000 428.200000 5.260000 429.280000 ;
      RECT 0.000000 427.760000 550.160000 428.200000 ;
      RECT 0.000000 426.780000 548.960000 427.760000 ;
      RECT 0.000000 426.560000 550.160000 426.780000 ;
      RECT 547.100000 425.480000 550.160000 426.560000 ;
      RECT 506.620000 425.480000 545.300000 426.560000 ;
      RECT 461.620000 425.480000 504.820000 426.560000 ;
      RECT 416.620000 425.480000 459.820000 426.560000 ;
      RECT 371.620000 425.480000 414.820000 426.560000 ;
      RECT 326.620000 425.480000 369.820000 426.560000 ;
      RECT 281.620000 425.480000 324.820000 426.560000 ;
      RECT 236.620000 425.480000 279.820000 426.560000 ;
      RECT 191.620000 425.480000 234.820000 426.560000 ;
      RECT 146.620000 425.480000 189.820000 426.560000 ;
      RECT 101.620000 425.480000 144.820000 426.560000 ;
      RECT 56.620000 425.480000 99.820000 426.560000 ;
      RECT 11.620000 425.480000 54.820000 426.560000 ;
      RECT 4.860000 425.480000 9.655000 426.560000 ;
      RECT 0.000000 425.480000 3.060000 426.560000 ;
      RECT 0.000000 424.100000 550.160000 425.480000 ;
      RECT 0.000000 423.840000 548.960000 424.100000 ;
      RECT 544.900000 423.120000 548.960000 423.840000 ;
      RECT 544.900000 422.760000 550.160000 423.120000 ;
      RECT 508.620000 422.760000 543.100000 423.840000 ;
      RECT 463.620000 422.760000 506.820000 423.840000 ;
      RECT 418.620000 422.760000 461.820000 423.840000 ;
      RECT 373.620000 422.760000 416.820000 423.840000 ;
      RECT 328.620000 422.760000 371.820000 423.840000 ;
      RECT 283.620000 422.760000 326.820000 423.840000 ;
      RECT 238.620000 422.760000 281.820000 423.840000 ;
      RECT 193.620000 422.760000 236.820000 423.840000 ;
      RECT 148.620000 422.760000 191.820000 423.840000 ;
      RECT 103.620000 422.760000 146.820000 423.840000 ;
      RECT 58.620000 422.760000 101.820000 423.840000 ;
      RECT 13.620000 422.760000 56.820000 423.840000 ;
      RECT 7.060000 422.760000 11.820000 423.840000 ;
      RECT 0.000000 422.760000 5.260000 423.840000 ;
      RECT 0.000000 421.120000 550.160000 422.760000 ;
      RECT 547.100000 420.440000 550.160000 421.120000 ;
      RECT 547.100000 420.040000 548.960000 420.440000 ;
      RECT 506.620000 420.040000 545.300000 421.120000 ;
      RECT 461.620000 420.040000 504.820000 421.120000 ;
      RECT 416.620000 420.040000 459.820000 421.120000 ;
      RECT 371.620000 420.040000 414.820000 421.120000 ;
      RECT 326.620000 420.040000 369.820000 421.120000 ;
      RECT 281.620000 420.040000 324.820000 421.120000 ;
      RECT 236.620000 420.040000 279.820000 421.120000 ;
      RECT 191.620000 420.040000 234.820000 421.120000 ;
      RECT 146.620000 420.040000 189.820000 421.120000 ;
      RECT 101.620000 420.040000 144.820000 421.120000 ;
      RECT 56.620000 420.040000 99.820000 421.120000 ;
      RECT 11.620000 420.040000 54.820000 421.120000 ;
      RECT 4.860000 420.040000 9.655000 421.120000 ;
      RECT 0.000000 420.040000 3.060000 421.120000 ;
      RECT 0.000000 419.460000 548.960000 420.040000 ;
      RECT 0.000000 418.400000 550.160000 419.460000 ;
      RECT 544.900000 417.390000 550.160000 418.400000 ;
      RECT 544.900000 417.320000 548.960000 417.390000 ;
      RECT 508.620000 417.320000 543.100000 418.400000 ;
      RECT 463.620000 417.320000 506.820000 418.400000 ;
      RECT 418.620000 417.320000 461.820000 418.400000 ;
      RECT 373.620000 417.320000 416.820000 418.400000 ;
      RECT 328.620000 417.320000 371.820000 418.400000 ;
      RECT 283.620000 417.320000 326.820000 418.400000 ;
      RECT 238.620000 417.320000 281.820000 418.400000 ;
      RECT 193.620000 417.320000 236.820000 418.400000 ;
      RECT 148.620000 417.320000 191.820000 418.400000 ;
      RECT 103.620000 417.320000 146.820000 418.400000 ;
      RECT 58.620000 417.320000 101.820000 418.400000 ;
      RECT 13.620000 417.320000 56.820000 418.400000 ;
      RECT 7.060000 417.320000 11.820000 418.400000 ;
      RECT 0.000000 417.320000 5.260000 418.400000 ;
      RECT 0.000000 416.410000 548.960000 417.320000 ;
      RECT 0.000000 415.680000 550.160000 416.410000 ;
      RECT 547.100000 414.600000 550.160000 415.680000 ;
      RECT 506.620000 414.600000 545.300000 415.680000 ;
      RECT 461.620000 414.600000 504.820000 415.680000 ;
      RECT 416.620000 414.600000 459.820000 415.680000 ;
      RECT 371.620000 414.600000 414.820000 415.680000 ;
      RECT 326.620000 414.600000 369.820000 415.680000 ;
      RECT 281.620000 414.600000 324.820000 415.680000 ;
      RECT 236.620000 414.600000 279.820000 415.680000 ;
      RECT 191.620000 414.600000 234.820000 415.680000 ;
      RECT 146.620000 414.600000 189.820000 415.680000 ;
      RECT 101.620000 414.600000 144.820000 415.680000 ;
      RECT 56.620000 414.600000 99.820000 415.680000 ;
      RECT 11.620000 414.600000 54.820000 415.680000 ;
      RECT 4.860000 414.600000 9.655000 415.680000 ;
      RECT 0.000000 414.600000 3.060000 415.680000 ;
      RECT 0.000000 413.730000 550.160000 414.600000 ;
      RECT 0.000000 412.960000 548.960000 413.730000 ;
      RECT 544.900000 412.750000 548.960000 412.960000 ;
      RECT 544.900000 411.880000 550.160000 412.750000 ;
      RECT 508.620000 411.880000 543.100000 412.960000 ;
      RECT 463.620000 411.880000 506.820000 412.960000 ;
      RECT 418.620000 411.880000 461.820000 412.960000 ;
      RECT 373.620000 411.880000 416.820000 412.960000 ;
      RECT 328.620000 411.880000 371.820000 412.960000 ;
      RECT 283.620000 411.880000 326.820000 412.960000 ;
      RECT 238.620000 411.880000 281.820000 412.960000 ;
      RECT 193.620000 411.880000 236.820000 412.960000 ;
      RECT 148.620000 411.880000 191.820000 412.960000 ;
      RECT 103.620000 411.880000 146.820000 412.960000 ;
      RECT 58.620000 411.880000 101.820000 412.960000 ;
      RECT 13.620000 411.880000 56.820000 412.960000 ;
      RECT 7.060000 411.880000 11.820000 412.960000 ;
      RECT 0.000000 411.880000 5.260000 412.960000 ;
      RECT 0.000000 410.240000 550.160000 411.880000 ;
      RECT 547.100000 410.070000 550.160000 410.240000 ;
      RECT 547.100000 409.160000 548.960000 410.070000 ;
      RECT 506.620000 409.160000 545.300000 410.240000 ;
      RECT 461.620000 409.160000 504.820000 410.240000 ;
      RECT 416.620000 409.160000 459.820000 410.240000 ;
      RECT 371.620000 409.160000 414.820000 410.240000 ;
      RECT 326.620000 409.160000 369.820000 410.240000 ;
      RECT 281.620000 409.160000 324.820000 410.240000 ;
      RECT 236.620000 409.160000 279.820000 410.240000 ;
      RECT 191.620000 409.160000 234.820000 410.240000 ;
      RECT 146.620000 409.160000 189.820000 410.240000 ;
      RECT 101.620000 409.160000 144.820000 410.240000 ;
      RECT 56.620000 409.160000 99.820000 410.240000 ;
      RECT 11.620000 409.160000 54.820000 410.240000 ;
      RECT 4.860000 409.160000 9.655000 410.240000 ;
      RECT 0.000000 409.160000 3.060000 410.240000 ;
      RECT 0.000000 409.090000 548.960000 409.160000 ;
      RECT 0.000000 407.520000 550.160000 409.090000 ;
      RECT 544.900000 407.020000 550.160000 407.520000 ;
      RECT 544.900000 406.440000 548.960000 407.020000 ;
      RECT 508.620000 406.440000 543.100000 407.520000 ;
      RECT 463.620000 406.440000 506.820000 407.520000 ;
      RECT 418.620000 406.440000 461.820000 407.520000 ;
      RECT 373.620000 406.440000 416.820000 407.520000 ;
      RECT 328.620000 406.440000 371.820000 407.520000 ;
      RECT 283.620000 406.440000 326.820000 407.520000 ;
      RECT 238.620000 406.440000 281.820000 407.520000 ;
      RECT 193.620000 406.440000 236.820000 407.520000 ;
      RECT 148.620000 406.440000 191.820000 407.520000 ;
      RECT 103.620000 406.440000 146.820000 407.520000 ;
      RECT 58.620000 406.440000 101.820000 407.520000 ;
      RECT 13.620000 406.440000 56.820000 407.520000 ;
      RECT 7.060000 406.440000 11.820000 407.520000 ;
      RECT 0.000000 406.440000 5.260000 407.520000 ;
      RECT 0.000000 406.040000 548.960000 406.440000 ;
      RECT 0.000000 404.800000 550.160000 406.040000 ;
      RECT 547.100000 403.720000 550.160000 404.800000 ;
      RECT 506.620000 403.720000 545.300000 404.800000 ;
      RECT 461.620000 403.720000 504.820000 404.800000 ;
      RECT 416.620000 403.720000 459.820000 404.800000 ;
      RECT 371.620000 403.720000 414.820000 404.800000 ;
      RECT 326.620000 403.720000 369.820000 404.800000 ;
      RECT 281.620000 403.720000 324.820000 404.800000 ;
      RECT 236.620000 403.720000 279.820000 404.800000 ;
      RECT 191.620000 403.720000 234.820000 404.800000 ;
      RECT 146.620000 403.720000 189.820000 404.800000 ;
      RECT 101.620000 403.720000 144.820000 404.800000 ;
      RECT 56.620000 403.720000 99.820000 404.800000 ;
      RECT 11.620000 403.720000 54.820000 404.800000 ;
      RECT 4.860000 403.720000 9.655000 404.800000 ;
      RECT 0.000000 403.720000 3.060000 404.800000 ;
      RECT 0.000000 403.360000 550.160000 403.720000 ;
      RECT 0.000000 402.380000 548.960000 403.360000 ;
      RECT 0.000000 402.080000 550.160000 402.380000 ;
      RECT 544.900000 401.000000 550.160000 402.080000 ;
      RECT 508.620000 401.000000 543.100000 402.080000 ;
      RECT 463.620000 401.000000 506.820000 402.080000 ;
      RECT 418.620000 401.000000 461.820000 402.080000 ;
      RECT 373.620000 401.000000 416.820000 402.080000 ;
      RECT 328.620000 401.000000 371.820000 402.080000 ;
      RECT 283.620000 401.000000 326.820000 402.080000 ;
      RECT 238.620000 401.000000 281.820000 402.080000 ;
      RECT 193.620000 401.000000 236.820000 402.080000 ;
      RECT 148.620000 401.000000 191.820000 402.080000 ;
      RECT 103.620000 401.000000 146.820000 402.080000 ;
      RECT 58.620000 401.000000 101.820000 402.080000 ;
      RECT 13.620000 401.000000 56.820000 402.080000 ;
      RECT 7.060000 401.000000 11.820000 402.080000 ;
      RECT 0.000000 401.000000 5.260000 402.080000 ;
      RECT 0.000000 399.700000 550.160000 401.000000 ;
      RECT 0.000000 399.360000 548.960000 399.700000 ;
      RECT 547.100000 398.720000 548.960000 399.360000 ;
      RECT 547.100000 398.280000 550.160000 398.720000 ;
      RECT 506.620000 398.280000 545.300000 399.360000 ;
      RECT 461.620000 398.280000 504.820000 399.360000 ;
      RECT 416.620000 398.280000 459.820000 399.360000 ;
      RECT 371.620000 398.280000 414.820000 399.360000 ;
      RECT 326.620000 398.280000 369.820000 399.360000 ;
      RECT 281.620000 398.280000 324.820000 399.360000 ;
      RECT 236.620000 398.280000 279.820000 399.360000 ;
      RECT 191.620000 398.280000 234.820000 399.360000 ;
      RECT 146.620000 398.280000 189.820000 399.360000 ;
      RECT 101.620000 398.280000 144.820000 399.360000 ;
      RECT 56.620000 398.280000 99.820000 399.360000 ;
      RECT 11.620000 398.280000 54.820000 399.360000 ;
      RECT 4.860000 398.280000 9.655000 399.360000 ;
      RECT 0.000000 398.280000 3.060000 399.360000 ;
      RECT 0.000000 396.650000 550.160000 398.280000 ;
      RECT 0.000000 396.640000 548.960000 396.650000 ;
      RECT 544.900000 395.670000 548.960000 396.640000 ;
      RECT 544.900000 395.560000 550.160000 395.670000 ;
      RECT 508.620000 395.560000 543.100000 396.640000 ;
      RECT 463.620000 395.560000 506.820000 396.640000 ;
      RECT 418.620000 395.560000 461.820000 396.640000 ;
      RECT 373.620000 395.560000 416.820000 396.640000 ;
      RECT 328.620000 395.560000 371.820000 396.640000 ;
      RECT 283.620000 395.560000 326.820000 396.640000 ;
      RECT 238.620000 395.560000 281.820000 396.640000 ;
      RECT 193.620000 395.560000 236.820000 396.640000 ;
      RECT 148.620000 395.560000 191.820000 396.640000 ;
      RECT 103.620000 395.560000 146.820000 396.640000 ;
      RECT 58.620000 395.560000 101.820000 396.640000 ;
      RECT 13.620000 395.560000 56.820000 396.640000 ;
      RECT 7.060000 395.560000 11.820000 396.640000 ;
      RECT 0.000000 395.560000 5.260000 396.640000 ;
      RECT 0.000000 393.920000 550.160000 395.560000 ;
      RECT 547.100000 392.990000 550.160000 393.920000 ;
      RECT 547.100000 392.840000 548.960000 392.990000 ;
      RECT 506.620000 392.840000 545.300000 393.920000 ;
      RECT 461.620000 392.840000 504.820000 393.920000 ;
      RECT 416.620000 392.840000 459.820000 393.920000 ;
      RECT 371.620000 392.840000 414.820000 393.920000 ;
      RECT 326.620000 392.840000 369.820000 393.920000 ;
      RECT 281.620000 392.840000 324.820000 393.920000 ;
      RECT 236.620000 392.840000 279.820000 393.920000 ;
      RECT 191.620000 392.840000 234.820000 393.920000 ;
      RECT 146.620000 392.840000 189.820000 393.920000 ;
      RECT 101.620000 392.840000 144.820000 393.920000 ;
      RECT 56.620000 392.840000 99.820000 393.920000 ;
      RECT 11.620000 392.840000 54.820000 393.920000 ;
      RECT 4.860000 392.840000 9.655000 393.920000 ;
      RECT 0.000000 392.840000 3.060000 393.920000 ;
      RECT 0.000000 392.010000 548.960000 392.840000 ;
      RECT 0.000000 391.200000 550.160000 392.010000 ;
      RECT 544.900000 390.120000 550.160000 391.200000 ;
      RECT 508.620000 390.120000 543.100000 391.200000 ;
      RECT 463.620000 390.120000 506.820000 391.200000 ;
      RECT 418.620000 390.120000 461.820000 391.200000 ;
      RECT 373.620000 390.120000 416.820000 391.200000 ;
      RECT 328.620000 390.120000 371.820000 391.200000 ;
      RECT 283.620000 390.120000 326.820000 391.200000 ;
      RECT 238.620000 390.120000 281.820000 391.200000 ;
      RECT 193.620000 390.120000 236.820000 391.200000 ;
      RECT 148.620000 390.120000 191.820000 391.200000 ;
      RECT 103.620000 390.120000 146.820000 391.200000 ;
      RECT 58.620000 390.120000 101.820000 391.200000 ;
      RECT 13.620000 390.120000 56.820000 391.200000 ;
      RECT 7.060000 390.120000 11.820000 391.200000 ;
      RECT 0.000000 390.120000 5.260000 391.200000 ;
      RECT 0.000000 389.940000 550.160000 390.120000 ;
      RECT 0.000000 388.960000 548.960000 389.940000 ;
      RECT 0.000000 388.480000 550.160000 388.960000 ;
      RECT 547.100000 387.400000 550.160000 388.480000 ;
      RECT 506.620000 387.400000 545.300000 388.480000 ;
      RECT 461.620000 387.400000 504.820000 388.480000 ;
      RECT 416.620000 387.400000 459.820000 388.480000 ;
      RECT 371.620000 387.400000 414.820000 388.480000 ;
      RECT 326.620000 387.400000 369.820000 388.480000 ;
      RECT 281.620000 387.400000 324.820000 388.480000 ;
      RECT 236.620000 387.400000 279.820000 388.480000 ;
      RECT 191.620000 387.400000 234.820000 388.480000 ;
      RECT 146.620000 387.400000 189.820000 388.480000 ;
      RECT 101.620000 387.400000 144.820000 388.480000 ;
      RECT 56.620000 387.400000 99.820000 388.480000 ;
      RECT 11.620000 387.400000 54.820000 388.480000 ;
      RECT 4.860000 387.400000 9.655000 388.480000 ;
      RECT 0.000000 387.400000 3.060000 388.480000 ;
      RECT 0.000000 386.280000 550.160000 387.400000 ;
      RECT 0.000000 385.760000 548.960000 386.280000 ;
      RECT 544.900000 385.300000 548.960000 385.760000 ;
      RECT 544.900000 384.680000 550.160000 385.300000 ;
      RECT 508.620000 384.680000 543.100000 385.760000 ;
      RECT 463.620000 384.680000 506.820000 385.760000 ;
      RECT 418.620000 384.680000 461.820000 385.760000 ;
      RECT 373.620000 384.680000 416.820000 385.760000 ;
      RECT 328.620000 384.680000 371.820000 385.760000 ;
      RECT 283.620000 384.680000 326.820000 385.760000 ;
      RECT 238.620000 384.680000 281.820000 385.760000 ;
      RECT 193.620000 384.680000 236.820000 385.760000 ;
      RECT 148.620000 384.680000 191.820000 385.760000 ;
      RECT 103.620000 384.680000 146.820000 385.760000 ;
      RECT 58.620000 384.680000 101.820000 385.760000 ;
      RECT 13.620000 384.680000 56.820000 385.760000 ;
      RECT 7.060000 384.680000 11.820000 385.760000 ;
      RECT 0.000000 384.680000 5.260000 385.760000 ;
      RECT 0.000000 383.040000 550.160000 384.680000 ;
      RECT 547.100000 382.620000 550.160000 383.040000 ;
      RECT 547.100000 381.960000 548.960000 382.620000 ;
      RECT 506.620000 381.960000 545.300000 383.040000 ;
      RECT 461.620000 381.960000 504.820000 383.040000 ;
      RECT 416.620000 381.960000 459.820000 383.040000 ;
      RECT 371.620000 381.960000 414.820000 383.040000 ;
      RECT 326.620000 381.960000 369.820000 383.040000 ;
      RECT 281.620000 381.960000 324.820000 383.040000 ;
      RECT 236.620000 381.960000 279.820000 383.040000 ;
      RECT 191.620000 381.960000 234.820000 383.040000 ;
      RECT 146.620000 381.960000 189.820000 383.040000 ;
      RECT 101.620000 381.960000 144.820000 383.040000 ;
      RECT 56.620000 381.960000 99.820000 383.040000 ;
      RECT 11.620000 381.960000 54.820000 383.040000 ;
      RECT 4.860000 381.960000 9.655000 383.040000 ;
      RECT 0.000000 381.960000 3.060000 383.040000 ;
      RECT 0.000000 381.640000 548.960000 381.960000 ;
      RECT 0.000000 380.320000 550.160000 381.640000 ;
      RECT 544.900000 379.570000 550.160000 380.320000 ;
      RECT 544.900000 379.240000 548.960000 379.570000 ;
      RECT 508.620000 379.240000 543.100000 380.320000 ;
      RECT 463.620000 379.240000 506.820000 380.320000 ;
      RECT 418.620000 379.240000 461.820000 380.320000 ;
      RECT 373.620000 379.240000 416.820000 380.320000 ;
      RECT 328.620000 379.240000 371.820000 380.320000 ;
      RECT 283.620000 379.240000 326.820000 380.320000 ;
      RECT 238.620000 379.240000 281.820000 380.320000 ;
      RECT 193.620000 379.240000 236.820000 380.320000 ;
      RECT 148.620000 379.240000 191.820000 380.320000 ;
      RECT 103.620000 379.240000 146.820000 380.320000 ;
      RECT 58.620000 379.240000 101.820000 380.320000 ;
      RECT 13.620000 379.240000 56.820000 380.320000 ;
      RECT 7.060000 379.240000 11.820000 380.320000 ;
      RECT 0.000000 379.240000 5.260000 380.320000 ;
      RECT 0.000000 378.590000 548.960000 379.240000 ;
      RECT 0.000000 377.600000 550.160000 378.590000 ;
      RECT 547.100000 376.520000 550.160000 377.600000 ;
      RECT 506.620000 376.520000 545.300000 377.600000 ;
      RECT 461.620000 376.520000 504.820000 377.600000 ;
      RECT 416.620000 376.520000 459.820000 377.600000 ;
      RECT 371.620000 376.520000 414.820000 377.600000 ;
      RECT 326.620000 376.520000 369.820000 377.600000 ;
      RECT 281.620000 376.520000 324.820000 377.600000 ;
      RECT 236.620000 376.520000 279.820000 377.600000 ;
      RECT 191.620000 376.520000 234.820000 377.600000 ;
      RECT 146.620000 376.520000 189.820000 377.600000 ;
      RECT 101.620000 376.520000 144.820000 377.600000 ;
      RECT 56.620000 376.520000 99.820000 377.600000 ;
      RECT 11.620000 376.520000 54.820000 377.600000 ;
      RECT 4.860000 376.520000 9.655000 377.600000 ;
      RECT 0.000000 376.520000 3.060000 377.600000 ;
      RECT 0.000000 375.910000 550.160000 376.520000 ;
      RECT 0.000000 374.930000 548.960000 375.910000 ;
      RECT 0.000000 374.880000 550.160000 374.930000 ;
      RECT 544.900000 373.800000 550.160000 374.880000 ;
      RECT 508.620000 373.800000 543.100000 374.880000 ;
      RECT 463.620000 373.800000 506.820000 374.880000 ;
      RECT 418.620000 373.800000 461.820000 374.880000 ;
      RECT 373.620000 373.800000 416.820000 374.880000 ;
      RECT 328.620000 373.800000 371.820000 374.880000 ;
      RECT 283.620000 373.800000 326.820000 374.880000 ;
      RECT 238.620000 373.800000 281.820000 374.880000 ;
      RECT 193.620000 373.800000 236.820000 374.880000 ;
      RECT 148.620000 373.800000 191.820000 374.880000 ;
      RECT 103.620000 373.800000 146.820000 374.880000 ;
      RECT 58.620000 373.800000 101.820000 374.880000 ;
      RECT 13.620000 373.800000 56.820000 374.880000 ;
      RECT 7.060000 373.800000 11.820000 374.880000 ;
      RECT 0.000000 373.800000 5.260000 374.880000 ;
      RECT 0.000000 372.250000 550.160000 373.800000 ;
      RECT 0.000000 372.160000 548.960000 372.250000 ;
      RECT 547.100000 371.270000 548.960000 372.160000 ;
      RECT 547.100000 371.080000 550.160000 371.270000 ;
      RECT 506.620000 371.080000 545.300000 372.160000 ;
      RECT 461.620000 371.080000 504.820000 372.160000 ;
      RECT 416.620000 371.080000 459.820000 372.160000 ;
      RECT 371.620000 371.080000 414.820000 372.160000 ;
      RECT 326.620000 371.080000 369.820000 372.160000 ;
      RECT 281.620000 371.080000 324.820000 372.160000 ;
      RECT 236.620000 371.080000 279.820000 372.160000 ;
      RECT 191.620000 371.080000 234.820000 372.160000 ;
      RECT 146.620000 371.080000 189.820000 372.160000 ;
      RECT 101.620000 371.080000 144.820000 372.160000 ;
      RECT 56.620000 371.080000 99.820000 372.160000 ;
      RECT 11.620000 371.080000 54.820000 372.160000 ;
      RECT 4.860000 371.080000 9.655000 372.160000 ;
      RECT 0.000000 371.080000 3.060000 372.160000 ;
      RECT 0.000000 369.440000 550.160000 371.080000 ;
      RECT 544.900000 369.200000 550.160000 369.440000 ;
      RECT 544.900000 368.360000 548.960000 369.200000 ;
      RECT 508.620000 368.360000 543.100000 369.440000 ;
      RECT 463.620000 368.360000 506.820000 369.440000 ;
      RECT 418.620000 368.360000 461.820000 369.440000 ;
      RECT 373.620000 368.360000 416.820000 369.440000 ;
      RECT 328.620000 368.360000 371.820000 369.440000 ;
      RECT 283.620000 368.360000 326.820000 369.440000 ;
      RECT 238.620000 368.360000 281.820000 369.440000 ;
      RECT 193.620000 368.360000 236.820000 369.440000 ;
      RECT 148.620000 368.360000 191.820000 369.440000 ;
      RECT 103.620000 368.360000 146.820000 369.440000 ;
      RECT 58.620000 368.360000 101.820000 369.440000 ;
      RECT 13.620000 368.360000 56.820000 369.440000 ;
      RECT 7.060000 368.360000 11.820000 369.440000 ;
      RECT 0.000000 368.360000 5.260000 369.440000 ;
      RECT 0.000000 368.220000 548.960000 368.360000 ;
      RECT 0.000000 366.720000 550.160000 368.220000 ;
      RECT 547.100000 365.640000 550.160000 366.720000 ;
      RECT 506.620000 365.640000 545.300000 366.720000 ;
      RECT 461.620000 365.640000 504.820000 366.720000 ;
      RECT 416.620000 365.640000 459.820000 366.720000 ;
      RECT 371.620000 365.640000 414.820000 366.720000 ;
      RECT 326.620000 365.640000 369.820000 366.720000 ;
      RECT 281.620000 365.640000 324.820000 366.720000 ;
      RECT 236.620000 365.640000 279.820000 366.720000 ;
      RECT 191.620000 365.640000 234.820000 366.720000 ;
      RECT 146.620000 365.640000 189.820000 366.720000 ;
      RECT 101.620000 365.640000 144.820000 366.720000 ;
      RECT 56.620000 365.640000 99.820000 366.720000 ;
      RECT 11.620000 365.640000 54.820000 366.720000 ;
      RECT 4.860000 365.640000 9.655000 366.720000 ;
      RECT 0.000000 365.640000 3.060000 366.720000 ;
      RECT 0.000000 365.540000 550.160000 365.640000 ;
      RECT 0.000000 364.560000 548.960000 365.540000 ;
      RECT 0.000000 364.000000 550.160000 364.560000 ;
      RECT 544.900000 362.920000 550.160000 364.000000 ;
      RECT 508.620000 362.920000 543.100000 364.000000 ;
      RECT 463.620000 362.920000 506.820000 364.000000 ;
      RECT 418.620000 362.920000 461.820000 364.000000 ;
      RECT 373.620000 362.920000 416.820000 364.000000 ;
      RECT 328.620000 362.920000 371.820000 364.000000 ;
      RECT 283.620000 362.920000 326.820000 364.000000 ;
      RECT 238.620000 362.920000 281.820000 364.000000 ;
      RECT 193.620000 362.920000 236.820000 364.000000 ;
      RECT 148.620000 362.920000 191.820000 364.000000 ;
      RECT 103.620000 362.920000 146.820000 364.000000 ;
      RECT 58.620000 362.920000 101.820000 364.000000 ;
      RECT 13.620000 362.920000 56.820000 364.000000 ;
      RECT 7.060000 362.920000 11.820000 364.000000 ;
      RECT 0.000000 362.920000 5.260000 364.000000 ;
      RECT 0.000000 361.880000 550.160000 362.920000 ;
      RECT 0.000000 361.280000 548.960000 361.880000 ;
      RECT 547.100000 360.900000 548.960000 361.280000 ;
      RECT 547.100000 360.200000 550.160000 360.900000 ;
      RECT 506.620000 360.200000 545.300000 361.280000 ;
      RECT 461.620000 360.200000 504.820000 361.280000 ;
      RECT 416.620000 360.200000 459.820000 361.280000 ;
      RECT 371.620000 360.200000 414.820000 361.280000 ;
      RECT 326.620000 360.200000 369.820000 361.280000 ;
      RECT 281.620000 360.200000 324.820000 361.280000 ;
      RECT 236.620000 360.200000 279.820000 361.280000 ;
      RECT 191.620000 360.200000 234.820000 361.280000 ;
      RECT 146.620000 360.200000 189.820000 361.280000 ;
      RECT 101.620000 360.200000 144.820000 361.280000 ;
      RECT 56.620000 360.200000 99.820000 361.280000 ;
      RECT 11.620000 360.200000 54.820000 361.280000 ;
      RECT 4.860000 360.200000 9.655000 361.280000 ;
      RECT 0.000000 360.200000 3.060000 361.280000 ;
      RECT 0.000000 358.830000 550.160000 360.200000 ;
      RECT 0.000000 358.560000 548.960000 358.830000 ;
      RECT 544.900000 357.850000 548.960000 358.560000 ;
      RECT 544.900000 357.480000 550.160000 357.850000 ;
      RECT 508.620000 357.480000 543.100000 358.560000 ;
      RECT 463.620000 357.480000 506.820000 358.560000 ;
      RECT 418.620000 357.480000 461.820000 358.560000 ;
      RECT 373.620000 357.480000 416.820000 358.560000 ;
      RECT 328.620000 357.480000 371.820000 358.560000 ;
      RECT 283.620000 357.480000 326.820000 358.560000 ;
      RECT 238.620000 357.480000 281.820000 358.560000 ;
      RECT 193.620000 357.480000 236.820000 358.560000 ;
      RECT 148.620000 357.480000 191.820000 358.560000 ;
      RECT 103.620000 357.480000 146.820000 358.560000 ;
      RECT 58.620000 357.480000 101.820000 358.560000 ;
      RECT 13.620000 357.480000 56.820000 358.560000 ;
      RECT 7.060000 357.480000 11.820000 358.560000 ;
      RECT 0.000000 357.480000 5.260000 358.560000 ;
      RECT 0.000000 355.840000 550.160000 357.480000 ;
      RECT 547.100000 355.170000 550.160000 355.840000 ;
      RECT 547.100000 354.760000 548.960000 355.170000 ;
      RECT 506.620000 354.760000 545.300000 355.840000 ;
      RECT 461.620000 354.760000 504.820000 355.840000 ;
      RECT 416.620000 354.760000 459.820000 355.840000 ;
      RECT 371.620000 354.760000 414.820000 355.840000 ;
      RECT 326.620000 354.760000 369.820000 355.840000 ;
      RECT 281.620000 354.760000 324.820000 355.840000 ;
      RECT 236.620000 354.760000 279.820000 355.840000 ;
      RECT 191.620000 354.760000 234.820000 355.840000 ;
      RECT 146.620000 354.760000 189.820000 355.840000 ;
      RECT 101.620000 354.760000 144.820000 355.840000 ;
      RECT 56.620000 354.760000 99.820000 355.840000 ;
      RECT 11.620000 354.760000 54.820000 355.840000 ;
      RECT 4.860000 354.760000 9.655000 355.840000 ;
      RECT 0.000000 354.760000 3.060000 355.840000 ;
      RECT 0.000000 354.190000 548.960000 354.760000 ;
      RECT 0.000000 353.120000 550.160000 354.190000 ;
      RECT 544.900000 352.040000 550.160000 353.120000 ;
      RECT 508.620000 352.040000 543.100000 353.120000 ;
      RECT 463.620000 352.040000 506.820000 353.120000 ;
      RECT 418.620000 352.040000 461.820000 353.120000 ;
      RECT 373.620000 352.040000 416.820000 353.120000 ;
      RECT 328.620000 352.040000 371.820000 353.120000 ;
      RECT 283.620000 352.040000 326.820000 353.120000 ;
      RECT 238.620000 352.040000 281.820000 353.120000 ;
      RECT 193.620000 352.040000 236.820000 353.120000 ;
      RECT 148.620000 352.040000 191.820000 353.120000 ;
      RECT 103.620000 352.040000 146.820000 353.120000 ;
      RECT 58.620000 352.040000 101.820000 353.120000 ;
      RECT 13.620000 352.040000 56.820000 353.120000 ;
      RECT 7.060000 352.040000 11.820000 353.120000 ;
      RECT 0.000000 352.040000 5.260000 353.120000 ;
      RECT 0.000000 351.510000 550.160000 352.040000 ;
      RECT 0.000000 350.530000 548.960000 351.510000 ;
      RECT 0.000000 350.400000 550.160000 350.530000 ;
      RECT 547.100000 349.320000 550.160000 350.400000 ;
      RECT 506.620000 349.320000 545.300000 350.400000 ;
      RECT 461.620000 349.320000 504.820000 350.400000 ;
      RECT 416.620000 349.320000 459.820000 350.400000 ;
      RECT 371.620000 349.320000 414.820000 350.400000 ;
      RECT 326.620000 349.320000 369.820000 350.400000 ;
      RECT 281.620000 349.320000 324.820000 350.400000 ;
      RECT 236.620000 349.320000 279.820000 350.400000 ;
      RECT 191.620000 349.320000 234.820000 350.400000 ;
      RECT 146.620000 349.320000 189.820000 350.400000 ;
      RECT 101.620000 349.320000 144.820000 350.400000 ;
      RECT 56.620000 349.320000 99.820000 350.400000 ;
      RECT 11.620000 349.320000 54.820000 350.400000 ;
      RECT 4.860000 349.320000 9.655000 350.400000 ;
      RECT 0.000000 349.320000 3.060000 350.400000 ;
      RECT 0.000000 348.460000 550.160000 349.320000 ;
      RECT 0.000000 347.680000 548.960000 348.460000 ;
      RECT 544.900000 347.480000 548.960000 347.680000 ;
      RECT 544.900000 346.600000 550.160000 347.480000 ;
      RECT 508.620000 346.600000 543.100000 347.680000 ;
      RECT 463.620000 346.600000 506.820000 347.680000 ;
      RECT 418.620000 346.600000 461.820000 347.680000 ;
      RECT 373.620000 346.600000 416.820000 347.680000 ;
      RECT 328.620000 346.600000 371.820000 347.680000 ;
      RECT 283.620000 346.600000 326.820000 347.680000 ;
      RECT 238.620000 346.600000 281.820000 347.680000 ;
      RECT 193.620000 346.600000 236.820000 347.680000 ;
      RECT 148.620000 346.600000 191.820000 347.680000 ;
      RECT 103.620000 346.600000 146.820000 347.680000 ;
      RECT 58.620000 346.600000 101.820000 347.680000 ;
      RECT 13.620000 346.600000 56.820000 347.680000 ;
      RECT 7.060000 346.600000 11.820000 347.680000 ;
      RECT 0.000000 346.600000 5.260000 347.680000 ;
      RECT 0.000000 344.960000 550.160000 346.600000 ;
      RECT 547.100000 344.800000 550.160000 344.960000 ;
      RECT 547.100000 343.880000 548.960000 344.800000 ;
      RECT 506.620000 343.880000 545.300000 344.960000 ;
      RECT 461.620000 343.880000 504.820000 344.960000 ;
      RECT 416.620000 343.880000 459.820000 344.960000 ;
      RECT 371.620000 343.880000 414.820000 344.960000 ;
      RECT 326.620000 343.880000 369.820000 344.960000 ;
      RECT 281.620000 343.880000 324.820000 344.960000 ;
      RECT 236.620000 343.880000 279.820000 344.960000 ;
      RECT 191.620000 343.880000 234.820000 344.960000 ;
      RECT 146.620000 343.880000 189.820000 344.960000 ;
      RECT 101.620000 343.880000 144.820000 344.960000 ;
      RECT 56.620000 343.880000 99.820000 344.960000 ;
      RECT 11.620000 343.880000 54.820000 344.960000 ;
      RECT 4.860000 343.880000 9.655000 344.960000 ;
      RECT 0.000000 343.880000 3.060000 344.960000 ;
      RECT 0.000000 343.820000 548.960000 343.880000 ;
      RECT 0.000000 342.240000 550.160000 343.820000 ;
      RECT 544.900000 341.160000 550.160000 342.240000 ;
      RECT 508.620000 341.160000 543.100000 342.240000 ;
      RECT 463.620000 341.160000 506.820000 342.240000 ;
      RECT 418.620000 341.160000 461.820000 342.240000 ;
      RECT 373.620000 341.160000 416.820000 342.240000 ;
      RECT 328.620000 341.160000 371.820000 342.240000 ;
      RECT 283.620000 341.160000 326.820000 342.240000 ;
      RECT 238.620000 341.160000 281.820000 342.240000 ;
      RECT 193.620000 341.160000 236.820000 342.240000 ;
      RECT 148.620000 341.160000 191.820000 342.240000 ;
      RECT 103.620000 341.160000 146.820000 342.240000 ;
      RECT 58.620000 341.160000 101.820000 342.240000 ;
      RECT 13.620000 341.160000 56.820000 342.240000 ;
      RECT 7.060000 341.160000 11.820000 342.240000 ;
      RECT 0.000000 341.160000 5.260000 342.240000 ;
      RECT 0.000000 341.140000 550.160000 341.160000 ;
      RECT 0.000000 340.160000 548.960000 341.140000 ;
      RECT 0.000000 339.520000 550.160000 340.160000 ;
      RECT 547.100000 338.440000 550.160000 339.520000 ;
      RECT 506.620000 338.440000 545.300000 339.520000 ;
      RECT 461.620000 338.440000 504.820000 339.520000 ;
      RECT 416.620000 338.440000 459.820000 339.520000 ;
      RECT 371.620000 338.440000 414.820000 339.520000 ;
      RECT 326.620000 338.440000 369.820000 339.520000 ;
      RECT 281.620000 338.440000 324.820000 339.520000 ;
      RECT 236.620000 338.440000 279.820000 339.520000 ;
      RECT 191.620000 338.440000 234.820000 339.520000 ;
      RECT 146.620000 338.440000 189.820000 339.520000 ;
      RECT 101.620000 338.440000 144.820000 339.520000 ;
      RECT 56.620000 338.440000 99.820000 339.520000 ;
      RECT 11.620000 338.440000 54.820000 339.520000 ;
      RECT 4.860000 338.440000 9.655000 339.520000 ;
      RECT 0.000000 338.440000 3.060000 339.520000 ;
      RECT 0.000000 338.090000 550.160000 338.440000 ;
      RECT 0.000000 337.110000 548.960000 338.090000 ;
      RECT 0.000000 336.800000 550.160000 337.110000 ;
      RECT 544.900000 335.720000 550.160000 336.800000 ;
      RECT 508.620000 335.720000 543.100000 336.800000 ;
      RECT 463.620000 335.720000 506.820000 336.800000 ;
      RECT 418.620000 335.720000 461.820000 336.800000 ;
      RECT 373.620000 335.720000 416.820000 336.800000 ;
      RECT 328.620000 335.720000 371.820000 336.800000 ;
      RECT 283.620000 335.720000 326.820000 336.800000 ;
      RECT 238.620000 335.720000 281.820000 336.800000 ;
      RECT 193.620000 335.720000 236.820000 336.800000 ;
      RECT 148.620000 335.720000 191.820000 336.800000 ;
      RECT 103.620000 335.720000 146.820000 336.800000 ;
      RECT 58.620000 335.720000 101.820000 336.800000 ;
      RECT 13.620000 335.720000 56.820000 336.800000 ;
      RECT 7.060000 335.720000 11.820000 336.800000 ;
      RECT 0.000000 335.720000 5.260000 336.800000 ;
      RECT 0.000000 334.430000 550.160000 335.720000 ;
      RECT 0.000000 334.080000 548.960000 334.430000 ;
      RECT 547.100000 333.450000 548.960000 334.080000 ;
      RECT 547.100000 333.000000 550.160000 333.450000 ;
      RECT 506.620000 333.000000 545.300000 334.080000 ;
      RECT 461.620000 333.000000 504.820000 334.080000 ;
      RECT 416.620000 333.000000 459.820000 334.080000 ;
      RECT 371.620000 333.000000 414.820000 334.080000 ;
      RECT 326.620000 333.000000 369.820000 334.080000 ;
      RECT 281.620000 333.000000 324.820000 334.080000 ;
      RECT 236.620000 333.000000 279.820000 334.080000 ;
      RECT 191.620000 333.000000 234.820000 334.080000 ;
      RECT 146.620000 333.000000 189.820000 334.080000 ;
      RECT 101.620000 333.000000 144.820000 334.080000 ;
      RECT 56.620000 333.000000 99.820000 334.080000 ;
      RECT 11.620000 333.000000 54.820000 334.080000 ;
      RECT 4.860000 333.000000 9.655000 334.080000 ;
      RECT 0.000000 333.000000 3.060000 334.080000 ;
      RECT 0.000000 331.360000 550.160000 333.000000 ;
      RECT 544.900000 330.770000 550.160000 331.360000 ;
      RECT 544.900000 330.280000 548.960000 330.770000 ;
      RECT 508.620000 330.280000 543.100000 331.360000 ;
      RECT 463.620000 330.280000 506.820000 331.360000 ;
      RECT 418.620000 330.280000 461.820000 331.360000 ;
      RECT 373.620000 330.280000 416.820000 331.360000 ;
      RECT 328.620000 330.280000 371.820000 331.360000 ;
      RECT 283.620000 330.280000 326.820000 331.360000 ;
      RECT 238.620000 330.280000 281.820000 331.360000 ;
      RECT 193.620000 330.280000 236.820000 331.360000 ;
      RECT 148.620000 330.280000 191.820000 331.360000 ;
      RECT 103.620000 330.280000 146.820000 331.360000 ;
      RECT 58.620000 330.280000 101.820000 331.360000 ;
      RECT 13.620000 330.280000 56.820000 331.360000 ;
      RECT 7.060000 330.280000 11.820000 331.360000 ;
      RECT 0.000000 330.280000 5.260000 331.360000 ;
      RECT 0.000000 329.790000 548.960000 330.280000 ;
      RECT 0.000000 328.640000 550.160000 329.790000 ;
      RECT 547.100000 327.720000 550.160000 328.640000 ;
      RECT 547.100000 327.560000 548.960000 327.720000 ;
      RECT 506.620000 327.560000 545.300000 328.640000 ;
      RECT 461.620000 327.560000 504.820000 328.640000 ;
      RECT 416.620000 327.560000 459.820000 328.640000 ;
      RECT 371.620000 327.560000 414.820000 328.640000 ;
      RECT 326.620000 327.560000 369.820000 328.640000 ;
      RECT 281.620000 327.560000 324.820000 328.640000 ;
      RECT 236.620000 327.560000 279.820000 328.640000 ;
      RECT 191.620000 327.560000 234.820000 328.640000 ;
      RECT 146.620000 327.560000 189.820000 328.640000 ;
      RECT 101.620000 327.560000 144.820000 328.640000 ;
      RECT 56.620000 327.560000 99.820000 328.640000 ;
      RECT 11.620000 327.560000 54.820000 328.640000 ;
      RECT 4.860000 327.560000 9.655000 328.640000 ;
      RECT 0.000000 327.560000 3.060000 328.640000 ;
      RECT 0.000000 326.740000 548.960000 327.560000 ;
      RECT 0.000000 325.920000 550.160000 326.740000 ;
      RECT 544.900000 324.840000 550.160000 325.920000 ;
      RECT 508.620000 324.840000 543.100000 325.920000 ;
      RECT 463.620000 324.840000 506.820000 325.920000 ;
      RECT 418.620000 324.840000 461.820000 325.920000 ;
      RECT 373.620000 324.840000 416.820000 325.920000 ;
      RECT 328.620000 324.840000 371.820000 325.920000 ;
      RECT 283.620000 324.840000 326.820000 325.920000 ;
      RECT 238.620000 324.840000 281.820000 325.920000 ;
      RECT 193.620000 324.840000 236.820000 325.920000 ;
      RECT 148.620000 324.840000 191.820000 325.920000 ;
      RECT 103.620000 324.840000 146.820000 325.920000 ;
      RECT 58.620000 324.840000 101.820000 325.920000 ;
      RECT 13.620000 324.840000 56.820000 325.920000 ;
      RECT 7.060000 324.840000 11.820000 325.920000 ;
      RECT 0.000000 324.840000 5.260000 325.920000 ;
      RECT 0.000000 324.060000 550.160000 324.840000 ;
      RECT 0.000000 323.200000 548.960000 324.060000 ;
      RECT 547.100000 323.080000 548.960000 323.200000 ;
      RECT 547.100000 322.120000 550.160000 323.080000 ;
      RECT 506.620000 322.120000 545.300000 323.200000 ;
      RECT 461.620000 322.120000 504.820000 323.200000 ;
      RECT 416.620000 322.120000 459.820000 323.200000 ;
      RECT 371.620000 322.120000 414.820000 323.200000 ;
      RECT 326.620000 322.120000 369.820000 323.200000 ;
      RECT 281.620000 322.120000 324.820000 323.200000 ;
      RECT 236.620000 322.120000 279.820000 323.200000 ;
      RECT 191.620000 322.120000 234.820000 323.200000 ;
      RECT 146.620000 322.120000 189.820000 323.200000 ;
      RECT 101.620000 322.120000 144.820000 323.200000 ;
      RECT 56.620000 322.120000 99.820000 323.200000 ;
      RECT 11.620000 322.120000 54.820000 323.200000 ;
      RECT 4.860000 322.120000 9.655000 323.200000 ;
      RECT 0.000000 322.120000 3.060000 323.200000 ;
      RECT 0.000000 320.480000 550.160000 322.120000 ;
      RECT 544.900000 320.400000 550.160000 320.480000 ;
      RECT 544.900000 319.420000 548.960000 320.400000 ;
      RECT 544.900000 319.400000 550.160000 319.420000 ;
      RECT 508.620000 319.400000 543.100000 320.480000 ;
      RECT 463.620000 319.400000 506.820000 320.480000 ;
      RECT 418.620000 319.400000 461.820000 320.480000 ;
      RECT 373.620000 319.400000 416.820000 320.480000 ;
      RECT 328.620000 319.400000 371.820000 320.480000 ;
      RECT 283.620000 319.400000 326.820000 320.480000 ;
      RECT 238.620000 319.400000 281.820000 320.480000 ;
      RECT 193.620000 319.400000 236.820000 320.480000 ;
      RECT 148.620000 319.400000 191.820000 320.480000 ;
      RECT 103.620000 319.400000 146.820000 320.480000 ;
      RECT 58.620000 319.400000 101.820000 320.480000 ;
      RECT 13.620000 319.400000 56.820000 320.480000 ;
      RECT 7.060000 319.400000 11.820000 320.480000 ;
      RECT 0.000000 319.400000 5.260000 320.480000 ;
      RECT 0.000000 317.760000 550.160000 319.400000 ;
      RECT 547.100000 317.350000 550.160000 317.760000 ;
      RECT 547.100000 316.680000 548.960000 317.350000 ;
      RECT 506.620000 316.680000 545.300000 317.760000 ;
      RECT 461.620000 316.680000 504.820000 317.760000 ;
      RECT 416.620000 316.680000 459.820000 317.760000 ;
      RECT 371.620000 316.680000 414.820000 317.760000 ;
      RECT 326.620000 316.680000 369.820000 317.760000 ;
      RECT 281.620000 316.680000 324.820000 317.760000 ;
      RECT 236.620000 316.680000 279.820000 317.760000 ;
      RECT 191.620000 316.680000 234.820000 317.760000 ;
      RECT 146.620000 316.680000 189.820000 317.760000 ;
      RECT 101.620000 316.680000 144.820000 317.760000 ;
      RECT 56.620000 316.680000 99.820000 317.760000 ;
      RECT 11.620000 316.680000 54.820000 317.760000 ;
      RECT 4.860000 316.680000 9.655000 317.760000 ;
      RECT 0.000000 316.680000 3.060000 317.760000 ;
      RECT 0.000000 316.370000 548.960000 316.680000 ;
      RECT 0.000000 315.040000 550.160000 316.370000 ;
      RECT 544.900000 313.960000 550.160000 315.040000 ;
      RECT 508.620000 313.960000 543.100000 315.040000 ;
      RECT 463.620000 313.960000 506.820000 315.040000 ;
      RECT 418.620000 313.960000 461.820000 315.040000 ;
      RECT 373.620000 313.960000 416.820000 315.040000 ;
      RECT 328.620000 313.960000 371.820000 315.040000 ;
      RECT 283.620000 313.960000 326.820000 315.040000 ;
      RECT 238.620000 313.960000 281.820000 315.040000 ;
      RECT 193.620000 313.960000 236.820000 315.040000 ;
      RECT 148.620000 313.960000 191.820000 315.040000 ;
      RECT 103.620000 313.960000 146.820000 315.040000 ;
      RECT 58.620000 313.960000 101.820000 315.040000 ;
      RECT 13.620000 313.960000 56.820000 315.040000 ;
      RECT 7.060000 313.960000 11.820000 315.040000 ;
      RECT 0.000000 313.960000 5.260000 315.040000 ;
      RECT 0.000000 313.690000 550.160000 313.960000 ;
      RECT 0.000000 312.710000 548.960000 313.690000 ;
      RECT 0.000000 312.320000 550.160000 312.710000 ;
      RECT 547.100000 311.240000 550.160000 312.320000 ;
      RECT 506.620000 311.240000 545.300000 312.320000 ;
      RECT 461.620000 311.240000 504.820000 312.320000 ;
      RECT 416.620000 311.240000 459.820000 312.320000 ;
      RECT 371.620000 311.240000 414.820000 312.320000 ;
      RECT 326.620000 311.240000 369.820000 312.320000 ;
      RECT 281.620000 311.240000 324.820000 312.320000 ;
      RECT 236.620000 311.240000 279.820000 312.320000 ;
      RECT 191.620000 311.240000 234.820000 312.320000 ;
      RECT 146.620000 311.240000 189.820000 312.320000 ;
      RECT 101.620000 311.240000 144.820000 312.320000 ;
      RECT 56.620000 311.240000 99.820000 312.320000 ;
      RECT 11.620000 311.240000 54.820000 312.320000 ;
      RECT 4.860000 311.240000 9.655000 312.320000 ;
      RECT 0.000000 311.240000 3.060000 312.320000 ;
      RECT 0.000000 310.030000 550.160000 311.240000 ;
      RECT 0.000000 309.600000 548.960000 310.030000 ;
      RECT 544.900000 309.050000 548.960000 309.600000 ;
      RECT 544.900000 308.520000 550.160000 309.050000 ;
      RECT 508.620000 308.520000 543.100000 309.600000 ;
      RECT 463.620000 308.520000 506.820000 309.600000 ;
      RECT 418.620000 308.520000 461.820000 309.600000 ;
      RECT 373.620000 308.520000 416.820000 309.600000 ;
      RECT 328.620000 308.520000 371.820000 309.600000 ;
      RECT 283.620000 308.520000 326.820000 309.600000 ;
      RECT 238.620000 308.520000 281.820000 309.600000 ;
      RECT 193.620000 308.520000 236.820000 309.600000 ;
      RECT 148.620000 308.520000 191.820000 309.600000 ;
      RECT 103.620000 308.520000 146.820000 309.600000 ;
      RECT 58.620000 308.520000 101.820000 309.600000 ;
      RECT 13.620000 308.520000 56.820000 309.600000 ;
      RECT 7.060000 308.520000 11.820000 309.600000 ;
      RECT 0.000000 308.520000 5.260000 309.600000 ;
      RECT 0.000000 306.980000 550.160000 308.520000 ;
      RECT 0.000000 306.880000 548.960000 306.980000 ;
      RECT 547.100000 306.000000 548.960000 306.880000 ;
      RECT 547.100000 305.800000 550.160000 306.000000 ;
      RECT 506.620000 305.800000 545.300000 306.880000 ;
      RECT 461.620000 305.800000 504.820000 306.880000 ;
      RECT 416.620000 305.800000 459.820000 306.880000 ;
      RECT 371.620000 305.800000 414.820000 306.880000 ;
      RECT 326.620000 305.800000 369.820000 306.880000 ;
      RECT 281.620000 305.800000 324.820000 306.880000 ;
      RECT 236.620000 305.800000 279.820000 306.880000 ;
      RECT 191.620000 305.800000 234.820000 306.880000 ;
      RECT 146.620000 305.800000 189.820000 306.880000 ;
      RECT 101.620000 305.800000 144.820000 306.880000 ;
      RECT 56.620000 305.800000 99.820000 306.880000 ;
      RECT 11.620000 305.800000 54.820000 306.880000 ;
      RECT 4.860000 305.800000 9.655000 306.880000 ;
      RECT 0.000000 305.800000 3.060000 306.880000 ;
      RECT 0.000000 304.160000 550.160000 305.800000 ;
      RECT 544.900000 303.320000 550.160000 304.160000 ;
      RECT 544.900000 303.080000 548.960000 303.320000 ;
      RECT 508.620000 303.080000 543.100000 304.160000 ;
      RECT 463.620000 303.080000 506.820000 304.160000 ;
      RECT 418.620000 303.080000 461.820000 304.160000 ;
      RECT 373.620000 303.080000 416.820000 304.160000 ;
      RECT 328.620000 303.080000 371.820000 304.160000 ;
      RECT 283.620000 303.080000 326.820000 304.160000 ;
      RECT 238.620000 303.080000 281.820000 304.160000 ;
      RECT 193.620000 303.080000 236.820000 304.160000 ;
      RECT 148.620000 303.080000 191.820000 304.160000 ;
      RECT 103.620000 303.080000 146.820000 304.160000 ;
      RECT 58.620000 303.080000 101.820000 304.160000 ;
      RECT 13.620000 303.080000 56.820000 304.160000 ;
      RECT 7.060000 303.080000 11.820000 304.160000 ;
      RECT 0.000000 303.080000 5.260000 304.160000 ;
      RECT 0.000000 302.340000 548.960000 303.080000 ;
      RECT 0.000000 301.440000 550.160000 302.340000 ;
      RECT 547.100000 300.360000 550.160000 301.440000 ;
      RECT 506.620000 300.360000 545.300000 301.440000 ;
      RECT 461.620000 300.360000 504.820000 301.440000 ;
      RECT 416.620000 300.360000 459.820000 301.440000 ;
      RECT 371.620000 300.360000 414.820000 301.440000 ;
      RECT 326.620000 300.360000 369.820000 301.440000 ;
      RECT 281.620000 300.360000 324.820000 301.440000 ;
      RECT 236.620000 300.360000 279.820000 301.440000 ;
      RECT 191.620000 300.360000 234.820000 301.440000 ;
      RECT 146.620000 300.360000 189.820000 301.440000 ;
      RECT 101.620000 300.360000 144.820000 301.440000 ;
      RECT 56.620000 300.360000 99.820000 301.440000 ;
      RECT 11.620000 300.360000 54.820000 301.440000 ;
      RECT 4.860000 300.360000 9.655000 301.440000 ;
      RECT 0.000000 300.360000 3.060000 301.440000 ;
      RECT 0.000000 300.270000 550.160000 300.360000 ;
      RECT 0.000000 299.290000 548.960000 300.270000 ;
      RECT 0.000000 298.720000 550.160000 299.290000 ;
      RECT 544.900000 297.640000 550.160000 298.720000 ;
      RECT 508.620000 297.640000 543.100000 298.720000 ;
      RECT 463.620000 297.640000 506.820000 298.720000 ;
      RECT 418.620000 297.640000 461.820000 298.720000 ;
      RECT 373.620000 297.640000 416.820000 298.720000 ;
      RECT 328.620000 297.640000 371.820000 298.720000 ;
      RECT 283.620000 297.640000 326.820000 298.720000 ;
      RECT 238.620000 297.640000 281.820000 298.720000 ;
      RECT 193.620000 297.640000 236.820000 298.720000 ;
      RECT 148.620000 297.640000 191.820000 298.720000 ;
      RECT 103.620000 297.640000 146.820000 298.720000 ;
      RECT 58.620000 297.640000 101.820000 298.720000 ;
      RECT 13.620000 297.640000 56.820000 298.720000 ;
      RECT 7.060000 297.640000 11.820000 298.720000 ;
      RECT 0.000000 297.640000 5.260000 298.720000 ;
      RECT 0.000000 296.610000 550.160000 297.640000 ;
      RECT 0.000000 296.000000 548.960000 296.610000 ;
      RECT 547.100000 295.630000 548.960000 296.000000 ;
      RECT 547.100000 294.920000 550.160000 295.630000 ;
      RECT 506.620000 294.920000 545.300000 296.000000 ;
      RECT 461.620000 294.920000 504.820000 296.000000 ;
      RECT 416.620000 294.920000 459.820000 296.000000 ;
      RECT 371.620000 294.920000 414.820000 296.000000 ;
      RECT 326.620000 294.920000 369.820000 296.000000 ;
      RECT 281.620000 294.920000 324.820000 296.000000 ;
      RECT 236.620000 294.920000 279.820000 296.000000 ;
      RECT 191.620000 294.920000 234.820000 296.000000 ;
      RECT 146.620000 294.920000 189.820000 296.000000 ;
      RECT 101.620000 294.920000 144.820000 296.000000 ;
      RECT 56.620000 294.920000 99.820000 296.000000 ;
      RECT 11.620000 294.920000 54.820000 296.000000 ;
      RECT 4.860000 294.920000 9.655000 296.000000 ;
      RECT 0.000000 294.920000 3.060000 296.000000 ;
      RECT 0.000000 293.280000 550.160000 294.920000 ;
      RECT 544.900000 292.950000 550.160000 293.280000 ;
      RECT 544.900000 292.200000 548.960000 292.950000 ;
      RECT 508.620000 292.200000 543.100000 293.280000 ;
      RECT 463.620000 292.200000 506.820000 293.280000 ;
      RECT 418.620000 292.200000 461.820000 293.280000 ;
      RECT 373.620000 292.200000 416.820000 293.280000 ;
      RECT 328.620000 292.200000 371.820000 293.280000 ;
      RECT 283.620000 292.200000 326.820000 293.280000 ;
      RECT 238.620000 292.200000 281.820000 293.280000 ;
      RECT 193.620000 292.200000 236.820000 293.280000 ;
      RECT 148.620000 292.200000 191.820000 293.280000 ;
      RECT 103.620000 292.200000 146.820000 293.280000 ;
      RECT 58.620000 292.200000 101.820000 293.280000 ;
      RECT 13.620000 292.200000 56.820000 293.280000 ;
      RECT 7.060000 292.200000 11.820000 293.280000 ;
      RECT 0.000000 292.200000 5.260000 293.280000 ;
      RECT 0.000000 291.970000 548.960000 292.200000 ;
      RECT 0.000000 290.560000 550.160000 291.970000 ;
      RECT 547.100000 289.900000 550.160000 290.560000 ;
      RECT 547.100000 289.480000 548.960000 289.900000 ;
      RECT 506.620000 289.480000 545.300000 290.560000 ;
      RECT 461.620000 289.480000 504.820000 290.560000 ;
      RECT 416.620000 289.480000 459.820000 290.560000 ;
      RECT 371.620000 289.480000 414.820000 290.560000 ;
      RECT 326.620000 289.480000 369.820000 290.560000 ;
      RECT 281.620000 289.480000 324.820000 290.560000 ;
      RECT 236.620000 289.480000 279.820000 290.560000 ;
      RECT 191.620000 289.480000 234.820000 290.560000 ;
      RECT 146.620000 289.480000 189.820000 290.560000 ;
      RECT 101.620000 289.480000 144.820000 290.560000 ;
      RECT 56.620000 289.480000 99.820000 290.560000 ;
      RECT 11.620000 289.480000 54.820000 290.560000 ;
      RECT 4.860000 289.480000 9.655000 290.560000 ;
      RECT 0.000000 289.480000 3.060000 290.560000 ;
      RECT 0.000000 288.920000 548.960000 289.480000 ;
      RECT 0.000000 287.840000 550.160000 288.920000 ;
      RECT 544.900000 286.760000 550.160000 287.840000 ;
      RECT 508.620000 286.760000 543.100000 287.840000 ;
      RECT 463.620000 286.760000 506.820000 287.840000 ;
      RECT 418.620000 286.760000 461.820000 287.840000 ;
      RECT 373.620000 286.760000 416.820000 287.840000 ;
      RECT 328.620000 286.760000 371.820000 287.840000 ;
      RECT 283.620000 286.760000 326.820000 287.840000 ;
      RECT 238.620000 286.760000 281.820000 287.840000 ;
      RECT 193.620000 286.760000 236.820000 287.840000 ;
      RECT 148.620000 286.760000 191.820000 287.840000 ;
      RECT 103.620000 286.760000 146.820000 287.840000 ;
      RECT 58.620000 286.760000 101.820000 287.840000 ;
      RECT 13.620000 286.760000 56.820000 287.840000 ;
      RECT 7.060000 286.760000 11.820000 287.840000 ;
      RECT 0.000000 286.760000 5.260000 287.840000 ;
      RECT 0.000000 286.240000 550.160000 286.760000 ;
      RECT 0.000000 285.260000 548.960000 286.240000 ;
      RECT 0.000000 285.120000 550.160000 285.260000 ;
      RECT 547.100000 284.040000 550.160000 285.120000 ;
      RECT 506.620000 284.040000 545.300000 285.120000 ;
      RECT 461.620000 284.040000 504.820000 285.120000 ;
      RECT 416.620000 284.040000 459.820000 285.120000 ;
      RECT 371.620000 284.040000 414.820000 285.120000 ;
      RECT 326.620000 284.040000 369.820000 285.120000 ;
      RECT 281.620000 284.040000 324.820000 285.120000 ;
      RECT 236.620000 284.040000 279.820000 285.120000 ;
      RECT 191.620000 284.040000 234.820000 285.120000 ;
      RECT 146.620000 284.040000 189.820000 285.120000 ;
      RECT 101.620000 284.040000 144.820000 285.120000 ;
      RECT 56.620000 284.040000 99.820000 285.120000 ;
      RECT 11.620000 284.040000 54.820000 285.120000 ;
      RECT 4.860000 284.040000 9.655000 285.120000 ;
      RECT 0.000000 284.040000 3.060000 285.120000 ;
      RECT 0.000000 282.580000 550.160000 284.040000 ;
      RECT 0.000000 282.400000 548.960000 282.580000 ;
      RECT 544.900000 281.600000 548.960000 282.400000 ;
      RECT 544.900000 281.320000 550.160000 281.600000 ;
      RECT 508.620000 281.320000 543.100000 282.400000 ;
      RECT 463.620000 281.320000 506.820000 282.400000 ;
      RECT 418.620000 281.320000 461.820000 282.400000 ;
      RECT 373.620000 281.320000 416.820000 282.400000 ;
      RECT 328.620000 281.320000 371.820000 282.400000 ;
      RECT 283.620000 281.320000 326.820000 282.400000 ;
      RECT 238.620000 281.320000 281.820000 282.400000 ;
      RECT 193.620000 281.320000 236.820000 282.400000 ;
      RECT 148.620000 281.320000 191.820000 282.400000 ;
      RECT 103.620000 281.320000 146.820000 282.400000 ;
      RECT 58.620000 281.320000 101.820000 282.400000 ;
      RECT 13.620000 281.320000 56.820000 282.400000 ;
      RECT 7.060000 281.320000 11.820000 282.400000 ;
      RECT 0.000000 281.320000 5.260000 282.400000 ;
      RECT 0.000000 279.680000 550.160000 281.320000 ;
      RECT 547.100000 279.530000 550.160000 279.680000 ;
      RECT 547.100000 278.600000 548.960000 279.530000 ;
      RECT 506.620000 278.600000 545.300000 279.680000 ;
      RECT 461.620000 278.600000 504.820000 279.680000 ;
      RECT 416.620000 278.600000 459.820000 279.680000 ;
      RECT 371.620000 278.600000 414.820000 279.680000 ;
      RECT 326.620000 278.600000 369.820000 279.680000 ;
      RECT 281.620000 278.600000 324.820000 279.680000 ;
      RECT 236.620000 278.600000 279.820000 279.680000 ;
      RECT 191.620000 278.600000 234.820000 279.680000 ;
      RECT 146.620000 278.600000 189.820000 279.680000 ;
      RECT 101.620000 278.600000 144.820000 279.680000 ;
      RECT 56.620000 278.600000 99.820000 279.680000 ;
      RECT 11.620000 278.600000 54.820000 279.680000 ;
      RECT 4.860000 278.600000 9.655000 279.680000 ;
      RECT 0.000000 278.600000 3.060000 279.680000 ;
      RECT 0.000000 278.550000 548.960000 278.600000 ;
      RECT 0.000000 276.960000 550.160000 278.550000 ;
      RECT 544.900000 275.880000 550.160000 276.960000 ;
      RECT 508.620000 275.880000 543.100000 276.960000 ;
      RECT 463.620000 275.880000 506.820000 276.960000 ;
      RECT 418.620000 275.880000 461.820000 276.960000 ;
      RECT 373.620000 275.880000 416.820000 276.960000 ;
      RECT 328.620000 275.880000 371.820000 276.960000 ;
      RECT 283.620000 275.880000 326.820000 276.960000 ;
      RECT 238.620000 275.880000 281.820000 276.960000 ;
      RECT 193.620000 275.880000 236.820000 276.960000 ;
      RECT 148.620000 275.880000 191.820000 276.960000 ;
      RECT 103.620000 275.880000 146.820000 276.960000 ;
      RECT 58.620000 275.880000 101.820000 276.960000 ;
      RECT 13.620000 275.880000 56.820000 276.960000 ;
      RECT 7.060000 275.880000 11.820000 276.960000 ;
      RECT 0.000000 275.880000 5.260000 276.960000 ;
      RECT 0.000000 275.870000 550.160000 275.880000 ;
      RECT 0.000000 274.890000 548.960000 275.870000 ;
      RECT 0.000000 274.240000 550.160000 274.890000 ;
      RECT 547.100000 273.160000 550.160000 274.240000 ;
      RECT 506.620000 273.160000 545.300000 274.240000 ;
      RECT 461.620000 273.160000 504.820000 274.240000 ;
      RECT 416.620000 273.160000 459.820000 274.240000 ;
      RECT 371.620000 273.160000 414.820000 274.240000 ;
      RECT 326.620000 273.160000 369.820000 274.240000 ;
      RECT 281.620000 273.160000 324.820000 274.240000 ;
      RECT 236.620000 273.160000 279.820000 274.240000 ;
      RECT 191.620000 273.160000 234.820000 274.240000 ;
      RECT 146.620000 273.160000 189.820000 274.240000 ;
      RECT 101.620000 273.160000 144.820000 274.240000 ;
      RECT 56.620000 273.160000 99.820000 274.240000 ;
      RECT 11.620000 273.160000 54.820000 274.240000 ;
      RECT 4.860000 273.160000 9.655000 274.240000 ;
      RECT 0.000000 273.160000 3.060000 274.240000 ;
      RECT 0.000000 272.210000 550.160000 273.160000 ;
      RECT 0.000000 271.520000 548.960000 272.210000 ;
      RECT 544.900000 271.230000 548.960000 271.520000 ;
      RECT 544.900000 270.440000 550.160000 271.230000 ;
      RECT 508.620000 270.440000 543.100000 271.520000 ;
      RECT 463.620000 270.440000 506.820000 271.520000 ;
      RECT 418.620000 270.440000 461.820000 271.520000 ;
      RECT 373.620000 270.440000 416.820000 271.520000 ;
      RECT 328.620000 270.440000 371.820000 271.520000 ;
      RECT 283.620000 270.440000 326.820000 271.520000 ;
      RECT 238.620000 270.440000 281.820000 271.520000 ;
      RECT 193.620000 270.440000 236.820000 271.520000 ;
      RECT 148.620000 270.440000 191.820000 271.520000 ;
      RECT 103.620000 270.440000 146.820000 271.520000 ;
      RECT 58.620000 270.440000 101.820000 271.520000 ;
      RECT 13.620000 270.440000 56.820000 271.520000 ;
      RECT 7.060000 270.440000 11.820000 271.520000 ;
      RECT 0.000000 270.440000 5.260000 271.520000 ;
      RECT 0.000000 269.160000 550.160000 270.440000 ;
      RECT 0.000000 268.800000 548.960000 269.160000 ;
      RECT 547.100000 268.180000 548.960000 268.800000 ;
      RECT 547.100000 267.720000 550.160000 268.180000 ;
      RECT 506.620000 267.720000 545.300000 268.800000 ;
      RECT 461.620000 267.720000 504.820000 268.800000 ;
      RECT 416.620000 267.720000 459.820000 268.800000 ;
      RECT 371.620000 267.720000 414.820000 268.800000 ;
      RECT 326.620000 267.720000 369.820000 268.800000 ;
      RECT 281.620000 267.720000 324.820000 268.800000 ;
      RECT 236.620000 267.720000 279.820000 268.800000 ;
      RECT 191.620000 267.720000 234.820000 268.800000 ;
      RECT 146.620000 267.720000 189.820000 268.800000 ;
      RECT 101.620000 267.720000 144.820000 268.800000 ;
      RECT 56.620000 267.720000 99.820000 268.800000 ;
      RECT 11.620000 267.720000 54.820000 268.800000 ;
      RECT 4.860000 267.720000 9.655000 268.800000 ;
      RECT 0.000000 267.720000 3.060000 268.800000 ;
      RECT 0.000000 266.080000 550.160000 267.720000 ;
      RECT 544.900000 265.500000 550.160000 266.080000 ;
      RECT 544.900000 265.000000 548.960000 265.500000 ;
      RECT 508.620000 265.000000 543.100000 266.080000 ;
      RECT 463.620000 265.000000 506.820000 266.080000 ;
      RECT 418.620000 265.000000 461.820000 266.080000 ;
      RECT 373.620000 265.000000 416.820000 266.080000 ;
      RECT 328.620000 265.000000 371.820000 266.080000 ;
      RECT 283.620000 265.000000 326.820000 266.080000 ;
      RECT 238.620000 265.000000 281.820000 266.080000 ;
      RECT 193.620000 265.000000 236.820000 266.080000 ;
      RECT 148.620000 265.000000 191.820000 266.080000 ;
      RECT 103.620000 265.000000 146.820000 266.080000 ;
      RECT 58.620000 265.000000 101.820000 266.080000 ;
      RECT 13.620000 265.000000 56.820000 266.080000 ;
      RECT 7.060000 265.000000 11.820000 266.080000 ;
      RECT 0.000000 265.000000 5.260000 266.080000 ;
      RECT 0.000000 264.520000 548.960000 265.000000 ;
      RECT 0.000000 263.360000 550.160000 264.520000 ;
      RECT 547.100000 262.280000 550.160000 263.360000 ;
      RECT 506.620000 262.280000 545.300000 263.360000 ;
      RECT 461.620000 262.280000 504.820000 263.360000 ;
      RECT 416.620000 262.280000 459.820000 263.360000 ;
      RECT 371.620000 262.280000 414.820000 263.360000 ;
      RECT 326.620000 262.280000 369.820000 263.360000 ;
      RECT 281.620000 262.280000 324.820000 263.360000 ;
      RECT 236.620000 262.280000 279.820000 263.360000 ;
      RECT 191.620000 262.280000 234.820000 263.360000 ;
      RECT 146.620000 262.280000 189.820000 263.360000 ;
      RECT 101.620000 262.280000 144.820000 263.360000 ;
      RECT 56.620000 262.280000 99.820000 263.360000 ;
      RECT 11.620000 262.280000 54.820000 263.360000 ;
      RECT 4.860000 262.280000 9.655000 263.360000 ;
      RECT 0.000000 262.280000 3.060000 263.360000 ;
      RECT 0.000000 261.840000 550.160000 262.280000 ;
      RECT 0.000000 260.860000 548.960000 261.840000 ;
      RECT 0.000000 260.640000 550.160000 260.860000 ;
      RECT 544.900000 259.560000 550.160000 260.640000 ;
      RECT 508.620000 259.560000 543.100000 260.640000 ;
      RECT 463.620000 259.560000 506.820000 260.640000 ;
      RECT 418.620000 259.560000 461.820000 260.640000 ;
      RECT 373.620000 259.560000 416.820000 260.640000 ;
      RECT 328.620000 259.560000 371.820000 260.640000 ;
      RECT 283.620000 259.560000 326.820000 260.640000 ;
      RECT 238.620000 259.560000 281.820000 260.640000 ;
      RECT 193.620000 259.560000 236.820000 260.640000 ;
      RECT 148.620000 259.560000 191.820000 260.640000 ;
      RECT 103.620000 259.560000 146.820000 260.640000 ;
      RECT 58.620000 259.560000 101.820000 260.640000 ;
      RECT 13.620000 259.560000 56.820000 260.640000 ;
      RECT 7.060000 259.560000 11.820000 260.640000 ;
      RECT 0.000000 259.560000 5.260000 260.640000 ;
      RECT 0.000000 258.790000 550.160000 259.560000 ;
      RECT 0.000000 257.920000 548.960000 258.790000 ;
      RECT 547.100000 257.810000 548.960000 257.920000 ;
      RECT 547.100000 256.840000 550.160000 257.810000 ;
      RECT 506.620000 256.840000 545.300000 257.920000 ;
      RECT 461.620000 256.840000 504.820000 257.920000 ;
      RECT 416.620000 256.840000 459.820000 257.920000 ;
      RECT 371.620000 256.840000 414.820000 257.920000 ;
      RECT 326.620000 256.840000 369.820000 257.920000 ;
      RECT 281.620000 256.840000 324.820000 257.920000 ;
      RECT 236.620000 256.840000 279.820000 257.920000 ;
      RECT 191.620000 256.840000 234.820000 257.920000 ;
      RECT 146.620000 256.840000 189.820000 257.920000 ;
      RECT 101.620000 256.840000 144.820000 257.920000 ;
      RECT 56.620000 256.840000 99.820000 257.920000 ;
      RECT 11.620000 256.840000 54.820000 257.920000 ;
      RECT 4.860000 256.840000 9.655000 257.920000 ;
      RECT 0.000000 256.840000 3.060000 257.920000 ;
      RECT 0.000000 255.200000 550.160000 256.840000 ;
      RECT 544.900000 255.130000 550.160000 255.200000 ;
      RECT 544.900000 254.150000 548.960000 255.130000 ;
      RECT 544.900000 254.120000 550.160000 254.150000 ;
      RECT 508.620000 254.120000 543.100000 255.200000 ;
      RECT 463.620000 254.120000 506.820000 255.200000 ;
      RECT 418.620000 254.120000 461.820000 255.200000 ;
      RECT 373.620000 254.120000 416.820000 255.200000 ;
      RECT 328.620000 254.120000 371.820000 255.200000 ;
      RECT 283.620000 254.120000 326.820000 255.200000 ;
      RECT 238.620000 254.120000 281.820000 255.200000 ;
      RECT 193.620000 254.120000 236.820000 255.200000 ;
      RECT 148.620000 254.120000 191.820000 255.200000 ;
      RECT 103.620000 254.120000 146.820000 255.200000 ;
      RECT 58.620000 254.120000 101.820000 255.200000 ;
      RECT 13.620000 254.120000 56.820000 255.200000 ;
      RECT 7.060000 254.120000 11.820000 255.200000 ;
      RECT 0.000000 254.120000 5.260000 255.200000 ;
      RECT 0.000000 252.480000 550.160000 254.120000 ;
      RECT 547.100000 251.470000 550.160000 252.480000 ;
      RECT 547.100000 251.400000 548.960000 251.470000 ;
      RECT 506.620000 251.400000 545.300000 252.480000 ;
      RECT 461.620000 251.400000 504.820000 252.480000 ;
      RECT 416.620000 251.400000 459.820000 252.480000 ;
      RECT 371.620000 251.400000 414.820000 252.480000 ;
      RECT 326.620000 251.400000 369.820000 252.480000 ;
      RECT 281.620000 251.400000 324.820000 252.480000 ;
      RECT 236.620000 251.400000 279.820000 252.480000 ;
      RECT 191.620000 251.400000 234.820000 252.480000 ;
      RECT 146.620000 251.400000 189.820000 252.480000 ;
      RECT 101.620000 251.400000 144.820000 252.480000 ;
      RECT 56.620000 251.400000 99.820000 252.480000 ;
      RECT 11.620000 251.400000 54.820000 252.480000 ;
      RECT 4.860000 251.400000 9.655000 252.480000 ;
      RECT 0.000000 251.400000 3.060000 252.480000 ;
      RECT 0.000000 250.490000 548.960000 251.400000 ;
      RECT 0.000000 249.760000 550.160000 250.490000 ;
      RECT 544.900000 248.680000 550.160000 249.760000 ;
      RECT 508.620000 248.680000 543.100000 249.760000 ;
      RECT 463.620000 248.680000 506.820000 249.760000 ;
      RECT 418.620000 248.680000 461.820000 249.760000 ;
      RECT 373.620000 248.680000 416.820000 249.760000 ;
      RECT 328.620000 248.680000 371.820000 249.760000 ;
      RECT 283.620000 248.680000 326.820000 249.760000 ;
      RECT 238.620000 248.680000 281.820000 249.760000 ;
      RECT 193.620000 248.680000 236.820000 249.760000 ;
      RECT 148.620000 248.680000 191.820000 249.760000 ;
      RECT 103.620000 248.680000 146.820000 249.760000 ;
      RECT 58.620000 248.680000 101.820000 249.760000 ;
      RECT 13.620000 248.680000 56.820000 249.760000 ;
      RECT 7.060000 248.680000 11.820000 249.760000 ;
      RECT 0.000000 248.680000 5.260000 249.760000 ;
      RECT 0.000000 248.420000 550.160000 248.680000 ;
      RECT 0.000000 247.440000 548.960000 248.420000 ;
      RECT 0.000000 247.040000 550.160000 247.440000 ;
      RECT 547.100000 245.960000 550.160000 247.040000 ;
      RECT 506.620000 245.960000 545.300000 247.040000 ;
      RECT 461.620000 245.960000 504.820000 247.040000 ;
      RECT 416.620000 245.960000 459.820000 247.040000 ;
      RECT 371.620000 245.960000 414.820000 247.040000 ;
      RECT 326.620000 245.960000 369.820000 247.040000 ;
      RECT 281.620000 245.960000 324.820000 247.040000 ;
      RECT 236.620000 245.960000 279.820000 247.040000 ;
      RECT 191.620000 245.960000 234.820000 247.040000 ;
      RECT 146.620000 245.960000 189.820000 247.040000 ;
      RECT 101.620000 245.960000 144.820000 247.040000 ;
      RECT 56.620000 245.960000 99.820000 247.040000 ;
      RECT 11.620000 245.960000 54.820000 247.040000 ;
      RECT 4.860000 245.960000 9.655000 247.040000 ;
      RECT 0.000000 245.960000 3.060000 247.040000 ;
      RECT 0.000000 244.760000 550.160000 245.960000 ;
      RECT 0.000000 244.320000 548.960000 244.760000 ;
      RECT 544.900000 243.780000 548.960000 244.320000 ;
      RECT 544.900000 243.240000 550.160000 243.780000 ;
      RECT 508.620000 243.240000 543.100000 244.320000 ;
      RECT 463.620000 243.240000 506.820000 244.320000 ;
      RECT 418.620000 243.240000 461.820000 244.320000 ;
      RECT 373.620000 243.240000 416.820000 244.320000 ;
      RECT 328.620000 243.240000 371.820000 244.320000 ;
      RECT 283.620000 243.240000 326.820000 244.320000 ;
      RECT 238.620000 243.240000 281.820000 244.320000 ;
      RECT 193.620000 243.240000 236.820000 244.320000 ;
      RECT 148.620000 243.240000 191.820000 244.320000 ;
      RECT 103.620000 243.240000 146.820000 244.320000 ;
      RECT 58.620000 243.240000 101.820000 244.320000 ;
      RECT 13.620000 243.240000 56.820000 244.320000 ;
      RECT 7.060000 243.240000 11.820000 244.320000 ;
      RECT 0.000000 243.240000 5.260000 244.320000 ;
      RECT 0.000000 241.600000 550.160000 243.240000 ;
      RECT 547.100000 241.100000 550.160000 241.600000 ;
      RECT 547.100000 240.520000 548.960000 241.100000 ;
      RECT 506.620000 240.520000 545.300000 241.600000 ;
      RECT 461.620000 240.520000 504.820000 241.600000 ;
      RECT 416.620000 240.520000 459.820000 241.600000 ;
      RECT 371.620000 240.520000 414.820000 241.600000 ;
      RECT 326.620000 240.520000 369.820000 241.600000 ;
      RECT 281.620000 240.520000 324.820000 241.600000 ;
      RECT 236.620000 240.520000 279.820000 241.600000 ;
      RECT 191.620000 240.520000 234.820000 241.600000 ;
      RECT 146.620000 240.520000 189.820000 241.600000 ;
      RECT 101.620000 240.520000 144.820000 241.600000 ;
      RECT 56.620000 240.520000 99.820000 241.600000 ;
      RECT 11.620000 240.520000 54.820000 241.600000 ;
      RECT 4.860000 240.520000 9.655000 241.600000 ;
      RECT 0.000000 240.520000 3.060000 241.600000 ;
      RECT 0.000000 240.120000 548.960000 240.520000 ;
      RECT 0.000000 238.880000 550.160000 240.120000 ;
      RECT 544.900000 238.050000 550.160000 238.880000 ;
      RECT 544.900000 237.800000 548.960000 238.050000 ;
      RECT 508.620000 237.800000 543.100000 238.880000 ;
      RECT 463.620000 237.800000 506.820000 238.880000 ;
      RECT 418.620000 237.800000 461.820000 238.880000 ;
      RECT 373.620000 237.800000 416.820000 238.880000 ;
      RECT 328.620000 237.800000 371.820000 238.880000 ;
      RECT 283.620000 237.800000 326.820000 238.880000 ;
      RECT 238.620000 237.800000 281.820000 238.880000 ;
      RECT 193.620000 237.800000 236.820000 238.880000 ;
      RECT 148.620000 237.800000 191.820000 238.880000 ;
      RECT 103.620000 237.800000 146.820000 238.880000 ;
      RECT 58.620000 237.800000 101.820000 238.880000 ;
      RECT 13.620000 237.800000 56.820000 238.880000 ;
      RECT 7.060000 237.800000 11.820000 238.880000 ;
      RECT 0.000000 237.800000 5.260000 238.880000 ;
      RECT 0.000000 237.070000 548.960000 237.800000 ;
      RECT 0.000000 236.160000 550.160000 237.070000 ;
      RECT 547.100000 235.080000 550.160000 236.160000 ;
      RECT 506.620000 235.080000 545.300000 236.160000 ;
      RECT 461.620000 235.080000 504.820000 236.160000 ;
      RECT 416.620000 235.080000 459.820000 236.160000 ;
      RECT 371.620000 235.080000 414.820000 236.160000 ;
      RECT 326.620000 235.080000 369.820000 236.160000 ;
      RECT 281.620000 235.080000 324.820000 236.160000 ;
      RECT 236.620000 235.080000 279.820000 236.160000 ;
      RECT 191.620000 235.080000 234.820000 236.160000 ;
      RECT 146.620000 235.080000 189.820000 236.160000 ;
      RECT 101.620000 235.080000 144.820000 236.160000 ;
      RECT 56.620000 235.080000 99.820000 236.160000 ;
      RECT 11.620000 235.080000 54.820000 236.160000 ;
      RECT 4.860000 235.080000 9.655000 236.160000 ;
      RECT 0.000000 235.080000 3.060000 236.160000 ;
      RECT 0.000000 234.390000 550.160000 235.080000 ;
      RECT 0.000000 233.440000 548.960000 234.390000 ;
      RECT 544.900000 233.410000 548.960000 233.440000 ;
      RECT 544.900000 232.360000 550.160000 233.410000 ;
      RECT 508.620000 232.360000 543.100000 233.440000 ;
      RECT 463.620000 232.360000 506.820000 233.440000 ;
      RECT 418.620000 232.360000 461.820000 233.440000 ;
      RECT 373.620000 232.360000 416.820000 233.440000 ;
      RECT 328.620000 232.360000 371.820000 233.440000 ;
      RECT 283.620000 232.360000 326.820000 233.440000 ;
      RECT 238.620000 232.360000 281.820000 233.440000 ;
      RECT 193.620000 232.360000 236.820000 233.440000 ;
      RECT 148.620000 232.360000 191.820000 233.440000 ;
      RECT 103.620000 232.360000 146.820000 233.440000 ;
      RECT 58.620000 232.360000 101.820000 233.440000 ;
      RECT 13.620000 232.360000 56.820000 233.440000 ;
      RECT 7.060000 232.360000 11.820000 233.440000 ;
      RECT 0.000000 232.360000 5.260000 233.440000 ;
      RECT 0.000000 230.730000 550.160000 232.360000 ;
      RECT 0.000000 230.720000 548.960000 230.730000 ;
      RECT 547.100000 229.750000 548.960000 230.720000 ;
      RECT 547.100000 229.640000 550.160000 229.750000 ;
      RECT 506.620000 229.640000 545.300000 230.720000 ;
      RECT 461.620000 229.640000 504.820000 230.720000 ;
      RECT 416.620000 229.640000 459.820000 230.720000 ;
      RECT 371.620000 229.640000 414.820000 230.720000 ;
      RECT 326.620000 229.640000 369.820000 230.720000 ;
      RECT 281.620000 229.640000 324.820000 230.720000 ;
      RECT 236.620000 229.640000 279.820000 230.720000 ;
      RECT 191.620000 229.640000 234.820000 230.720000 ;
      RECT 146.620000 229.640000 189.820000 230.720000 ;
      RECT 101.620000 229.640000 144.820000 230.720000 ;
      RECT 56.620000 229.640000 99.820000 230.720000 ;
      RECT 11.620000 229.640000 54.820000 230.720000 ;
      RECT 4.860000 229.640000 9.655000 230.720000 ;
      RECT 0.000000 229.640000 3.060000 230.720000 ;
      RECT 0.000000 228.000000 550.160000 229.640000 ;
      RECT 544.900000 227.680000 550.160000 228.000000 ;
      RECT 544.900000 226.920000 548.960000 227.680000 ;
      RECT 508.620000 226.920000 543.100000 228.000000 ;
      RECT 463.620000 226.920000 506.820000 228.000000 ;
      RECT 418.620000 226.920000 461.820000 228.000000 ;
      RECT 373.620000 226.920000 416.820000 228.000000 ;
      RECT 328.620000 226.920000 371.820000 228.000000 ;
      RECT 283.620000 226.920000 326.820000 228.000000 ;
      RECT 238.620000 226.920000 281.820000 228.000000 ;
      RECT 193.620000 226.920000 236.820000 228.000000 ;
      RECT 148.620000 226.920000 191.820000 228.000000 ;
      RECT 103.620000 226.920000 146.820000 228.000000 ;
      RECT 58.620000 226.920000 101.820000 228.000000 ;
      RECT 13.620000 226.920000 56.820000 228.000000 ;
      RECT 7.060000 226.920000 11.820000 228.000000 ;
      RECT 0.000000 226.920000 5.260000 228.000000 ;
      RECT 0.000000 226.700000 548.960000 226.920000 ;
      RECT 0.000000 225.280000 550.160000 226.700000 ;
      RECT 547.100000 224.200000 550.160000 225.280000 ;
      RECT 506.620000 224.200000 545.300000 225.280000 ;
      RECT 461.620000 224.200000 504.820000 225.280000 ;
      RECT 416.620000 224.200000 459.820000 225.280000 ;
      RECT 371.620000 224.200000 414.820000 225.280000 ;
      RECT 326.620000 224.200000 369.820000 225.280000 ;
      RECT 281.620000 224.200000 324.820000 225.280000 ;
      RECT 236.620000 224.200000 279.820000 225.280000 ;
      RECT 191.620000 224.200000 234.820000 225.280000 ;
      RECT 146.620000 224.200000 189.820000 225.280000 ;
      RECT 101.620000 224.200000 144.820000 225.280000 ;
      RECT 56.620000 224.200000 99.820000 225.280000 ;
      RECT 11.620000 224.200000 54.820000 225.280000 ;
      RECT 4.860000 224.200000 9.655000 225.280000 ;
      RECT 0.000000 224.200000 3.060000 225.280000 ;
      RECT 0.000000 224.020000 550.160000 224.200000 ;
      RECT 0.000000 223.040000 548.960000 224.020000 ;
      RECT 0.000000 222.560000 550.160000 223.040000 ;
      RECT 544.900000 221.480000 550.160000 222.560000 ;
      RECT 508.620000 221.480000 543.100000 222.560000 ;
      RECT 463.620000 221.480000 506.820000 222.560000 ;
      RECT 418.620000 221.480000 461.820000 222.560000 ;
      RECT 373.620000 221.480000 416.820000 222.560000 ;
      RECT 328.620000 221.480000 371.820000 222.560000 ;
      RECT 283.620000 221.480000 326.820000 222.560000 ;
      RECT 238.620000 221.480000 281.820000 222.560000 ;
      RECT 193.620000 221.480000 236.820000 222.560000 ;
      RECT 148.620000 221.480000 191.820000 222.560000 ;
      RECT 103.620000 221.480000 146.820000 222.560000 ;
      RECT 58.620000 221.480000 101.820000 222.560000 ;
      RECT 13.620000 221.480000 56.820000 222.560000 ;
      RECT 7.060000 221.480000 11.820000 222.560000 ;
      RECT 0.000000 221.480000 5.260000 222.560000 ;
      RECT 0.000000 220.360000 550.160000 221.480000 ;
      RECT 0.000000 219.840000 548.960000 220.360000 ;
      RECT 547.100000 219.380000 548.960000 219.840000 ;
      RECT 547.100000 218.760000 550.160000 219.380000 ;
      RECT 506.620000 218.760000 545.300000 219.840000 ;
      RECT 461.620000 218.760000 504.820000 219.840000 ;
      RECT 416.620000 218.760000 459.820000 219.840000 ;
      RECT 371.620000 218.760000 414.820000 219.840000 ;
      RECT 326.620000 218.760000 369.820000 219.840000 ;
      RECT 281.620000 218.760000 324.820000 219.840000 ;
      RECT 236.620000 218.760000 279.820000 219.840000 ;
      RECT 191.620000 218.760000 234.820000 219.840000 ;
      RECT 146.620000 218.760000 189.820000 219.840000 ;
      RECT 101.620000 218.760000 144.820000 219.840000 ;
      RECT 56.620000 218.760000 99.820000 219.840000 ;
      RECT 11.620000 218.760000 54.820000 219.840000 ;
      RECT 4.860000 218.760000 9.655000 219.840000 ;
      RECT 0.000000 218.760000 3.060000 219.840000 ;
      RECT 0.000000 217.310000 550.160000 218.760000 ;
      RECT 0.000000 217.120000 548.960000 217.310000 ;
      RECT 544.900000 216.330000 548.960000 217.120000 ;
      RECT 544.900000 216.040000 550.160000 216.330000 ;
      RECT 508.620000 216.040000 543.100000 217.120000 ;
      RECT 463.620000 216.040000 506.820000 217.120000 ;
      RECT 418.620000 216.040000 461.820000 217.120000 ;
      RECT 373.620000 216.040000 416.820000 217.120000 ;
      RECT 328.620000 216.040000 371.820000 217.120000 ;
      RECT 283.620000 216.040000 326.820000 217.120000 ;
      RECT 238.620000 216.040000 281.820000 217.120000 ;
      RECT 193.620000 216.040000 236.820000 217.120000 ;
      RECT 148.620000 216.040000 191.820000 217.120000 ;
      RECT 103.620000 216.040000 146.820000 217.120000 ;
      RECT 58.620000 216.040000 101.820000 217.120000 ;
      RECT 13.620000 216.040000 56.820000 217.120000 ;
      RECT 7.060000 216.040000 11.820000 217.120000 ;
      RECT 0.000000 216.040000 5.260000 217.120000 ;
      RECT 0.000000 214.400000 550.160000 216.040000 ;
      RECT 547.100000 213.650000 550.160000 214.400000 ;
      RECT 547.100000 213.320000 548.960000 213.650000 ;
      RECT 506.620000 213.320000 545.300000 214.400000 ;
      RECT 461.620000 213.320000 504.820000 214.400000 ;
      RECT 416.620000 213.320000 459.820000 214.400000 ;
      RECT 371.620000 213.320000 414.820000 214.400000 ;
      RECT 326.620000 213.320000 369.820000 214.400000 ;
      RECT 281.620000 213.320000 324.820000 214.400000 ;
      RECT 236.620000 213.320000 279.820000 214.400000 ;
      RECT 191.620000 213.320000 234.820000 214.400000 ;
      RECT 146.620000 213.320000 189.820000 214.400000 ;
      RECT 101.620000 213.320000 144.820000 214.400000 ;
      RECT 56.620000 213.320000 99.820000 214.400000 ;
      RECT 11.620000 213.320000 54.820000 214.400000 ;
      RECT 4.860000 213.320000 9.655000 214.400000 ;
      RECT 0.000000 213.320000 3.060000 214.400000 ;
      RECT 0.000000 212.670000 548.960000 213.320000 ;
      RECT 0.000000 211.680000 550.160000 212.670000 ;
      RECT 544.900000 210.600000 550.160000 211.680000 ;
      RECT 508.620000 210.600000 543.100000 211.680000 ;
      RECT 463.620000 210.600000 506.820000 211.680000 ;
      RECT 418.620000 210.600000 461.820000 211.680000 ;
      RECT 373.620000 210.600000 416.820000 211.680000 ;
      RECT 328.620000 210.600000 371.820000 211.680000 ;
      RECT 283.620000 210.600000 326.820000 211.680000 ;
      RECT 238.620000 210.600000 281.820000 211.680000 ;
      RECT 193.620000 210.600000 236.820000 211.680000 ;
      RECT 148.620000 210.600000 191.820000 211.680000 ;
      RECT 103.620000 210.600000 146.820000 211.680000 ;
      RECT 58.620000 210.600000 101.820000 211.680000 ;
      RECT 13.620000 210.600000 56.820000 211.680000 ;
      RECT 7.060000 210.600000 11.820000 211.680000 ;
      RECT 0.000000 210.600000 5.260000 211.680000 ;
      RECT 0.000000 209.990000 550.160000 210.600000 ;
      RECT 0.000000 209.010000 548.960000 209.990000 ;
      RECT 0.000000 208.960000 550.160000 209.010000 ;
      RECT 547.100000 207.880000 550.160000 208.960000 ;
      RECT 506.620000 207.880000 545.300000 208.960000 ;
      RECT 461.620000 207.880000 504.820000 208.960000 ;
      RECT 416.620000 207.880000 459.820000 208.960000 ;
      RECT 371.620000 207.880000 414.820000 208.960000 ;
      RECT 326.620000 207.880000 369.820000 208.960000 ;
      RECT 281.620000 207.880000 324.820000 208.960000 ;
      RECT 236.620000 207.880000 279.820000 208.960000 ;
      RECT 191.620000 207.880000 234.820000 208.960000 ;
      RECT 146.620000 207.880000 189.820000 208.960000 ;
      RECT 101.620000 207.880000 144.820000 208.960000 ;
      RECT 56.620000 207.880000 99.820000 208.960000 ;
      RECT 11.620000 207.880000 54.820000 208.960000 ;
      RECT 4.860000 207.880000 9.655000 208.960000 ;
      RECT 0.000000 207.880000 3.060000 208.960000 ;
      RECT 0.000000 206.940000 550.160000 207.880000 ;
      RECT 0.000000 206.240000 548.960000 206.940000 ;
      RECT 544.900000 205.960000 548.960000 206.240000 ;
      RECT 544.900000 205.160000 550.160000 205.960000 ;
      RECT 508.620000 205.160000 543.100000 206.240000 ;
      RECT 463.620000 205.160000 506.820000 206.240000 ;
      RECT 418.620000 205.160000 461.820000 206.240000 ;
      RECT 373.620000 205.160000 416.820000 206.240000 ;
      RECT 328.620000 205.160000 371.820000 206.240000 ;
      RECT 283.620000 205.160000 326.820000 206.240000 ;
      RECT 238.620000 205.160000 281.820000 206.240000 ;
      RECT 193.620000 205.160000 236.820000 206.240000 ;
      RECT 148.620000 205.160000 191.820000 206.240000 ;
      RECT 103.620000 205.160000 146.820000 206.240000 ;
      RECT 58.620000 205.160000 101.820000 206.240000 ;
      RECT 13.620000 205.160000 56.820000 206.240000 ;
      RECT 7.060000 205.160000 11.820000 206.240000 ;
      RECT 0.000000 205.160000 5.260000 206.240000 ;
      RECT 0.000000 203.520000 550.160000 205.160000 ;
      RECT 547.100000 203.280000 550.160000 203.520000 ;
      RECT 547.100000 202.440000 548.960000 203.280000 ;
      RECT 506.620000 202.440000 545.300000 203.520000 ;
      RECT 461.620000 202.440000 504.820000 203.520000 ;
      RECT 416.620000 202.440000 459.820000 203.520000 ;
      RECT 371.620000 202.440000 414.820000 203.520000 ;
      RECT 326.620000 202.440000 369.820000 203.520000 ;
      RECT 281.620000 202.440000 324.820000 203.520000 ;
      RECT 236.620000 202.440000 279.820000 203.520000 ;
      RECT 191.620000 202.440000 234.820000 203.520000 ;
      RECT 146.620000 202.440000 189.820000 203.520000 ;
      RECT 101.620000 202.440000 144.820000 203.520000 ;
      RECT 56.620000 202.440000 99.820000 203.520000 ;
      RECT 11.620000 202.440000 54.820000 203.520000 ;
      RECT 4.860000 202.440000 9.655000 203.520000 ;
      RECT 0.000000 202.440000 3.060000 203.520000 ;
      RECT 0.000000 202.300000 548.960000 202.440000 ;
      RECT 0.000000 200.800000 550.160000 202.300000 ;
      RECT 544.900000 200.230000 550.160000 200.800000 ;
      RECT 544.900000 199.720000 548.960000 200.230000 ;
      RECT 508.620000 199.720000 543.100000 200.800000 ;
      RECT 463.620000 199.720000 506.820000 200.800000 ;
      RECT 418.620000 199.720000 461.820000 200.800000 ;
      RECT 373.620000 199.720000 416.820000 200.800000 ;
      RECT 328.620000 199.720000 371.820000 200.800000 ;
      RECT 283.620000 199.720000 326.820000 200.800000 ;
      RECT 238.620000 199.720000 281.820000 200.800000 ;
      RECT 193.620000 199.720000 236.820000 200.800000 ;
      RECT 148.620000 199.720000 191.820000 200.800000 ;
      RECT 103.620000 199.720000 146.820000 200.800000 ;
      RECT 58.620000 199.720000 101.820000 200.800000 ;
      RECT 13.620000 199.720000 56.820000 200.800000 ;
      RECT 7.060000 199.720000 11.820000 200.800000 ;
      RECT 0.000000 199.720000 5.260000 200.800000 ;
      RECT 0.000000 199.250000 548.960000 199.720000 ;
      RECT 0.000000 198.080000 550.160000 199.250000 ;
      RECT 547.100000 197.000000 550.160000 198.080000 ;
      RECT 506.620000 197.000000 545.300000 198.080000 ;
      RECT 461.620000 197.000000 504.820000 198.080000 ;
      RECT 416.620000 197.000000 459.820000 198.080000 ;
      RECT 371.620000 197.000000 414.820000 198.080000 ;
      RECT 326.620000 197.000000 369.820000 198.080000 ;
      RECT 281.620000 197.000000 324.820000 198.080000 ;
      RECT 236.620000 197.000000 279.820000 198.080000 ;
      RECT 191.620000 197.000000 234.820000 198.080000 ;
      RECT 146.620000 197.000000 189.820000 198.080000 ;
      RECT 101.620000 197.000000 144.820000 198.080000 ;
      RECT 56.620000 197.000000 99.820000 198.080000 ;
      RECT 11.620000 197.000000 54.820000 198.080000 ;
      RECT 4.860000 197.000000 9.655000 198.080000 ;
      RECT 0.000000 197.000000 3.060000 198.080000 ;
      RECT 0.000000 196.570000 550.160000 197.000000 ;
      RECT 0.000000 195.590000 548.960000 196.570000 ;
      RECT 0.000000 195.360000 550.160000 195.590000 ;
      RECT 544.900000 194.280000 550.160000 195.360000 ;
      RECT 508.620000 194.280000 543.100000 195.360000 ;
      RECT 463.620000 194.280000 506.820000 195.360000 ;
      RECT 418.620000 194.280000 461.820000 195.360000 ;
      RECT 373.620000 194.280000 416.820000 195.360000 ;
      RECT 328.620000 194.280000 371.820000 195.360000 ;
      RECT 283.620000 194.280000 326.820000 195.360000 ;
      RECT 238.620000 194.280000 281.820000 195.360000 ;
      RECT 193.620000 194.280000 236.820000 195.360000 ;
      RECT 148.620000 194.280000 191.820000 195.360000 ;
      RECT 103.620000 194.280000 146.820000 195.360000 ;
      RECT 58.620000 194.280000 101.820000 195.360000 ;
      RECT 13.620000 194.280000 56.820000 195.360000 ;
      RECT 7.060000 194.280000 11.820000 195.360000 ;
      RECT 0.000000 194.280000 5.260000 195.360000 ;
      RECT 0.000000 192.910000 550.160000 194.280000 ;
      RECT 0.000000 192.640000 548.960000 192.910000 ;
      RECT 547.100000 191.930000 548.960000 192.640000 ;
      RECT 547.100000 191.560000 550.160000 191.930000 ;
      RECT 506.620000 191.560000 545.300000 192.640000 ;
      RECT 461.620000 191.560000 504.820000 192.640000 ;
      RECT 416.620000 191.560000 459.820000 192.640000 ;
      RECT 371.620000 191.560000 414.820000 192.640000 ;
      RECT 326.620000 191.560000 369.820000 192.640000 ;
      RECT 281.620000 191.560000 324.820000 192.640000 ;
      RECT 236.620000 191.560000 279.820000 192.640000 ;
      RECT 191.620000 191.560000 234.820000 192.640000 ;
      RECT 146.620000 191.560000 189.820000 192.640000 ;
      RECT 101.620000 191.560000 144.820000 192.640000 ;
      RECT 56.620000 191.560000 99.820000 192.640000 ;
      RECT 11.620000 191.560000 54.820000 192.640000 ;
      RECT 4.860000 191.560000 9.655000 192.640000 ;
      RECT 0.000000 191.560000 3.060000 192.640000 ;
      RECT 0.000000 189.920000 550.160000 191.560000 ;
      RECT 544.900000 189.860000 550.160000 189.920000 ;
      RECT 544.900000 188.880000 548.960000 189.860000 ;
      RECT 544.900000 188.840000 550.160000 188.880000 ;
      RECT 508.620000 188.840000 543.100000 189.920000 ;
      RECT 463.620000 188.840000 506.820000 189.920000 ;
      RECT 418.620000 188.840000 461.820000 189.920000 ;
      RECT 373.620000 188.840000 416.820000 189.920000 ;
      RECT 328.620000 188.840000 371.820000 189.920000 ;
      RECT 283.620000 188.840000 326.820000 189.920000 ;
      RECT 238.620000 188.840000 281.820000 189.920000 ;
      RECT 193.620000 188.840000 236.820000 189.920000 ;
      RECT 148.620000 188.840000 191.820000 189.920000 ;
      RECT 103.620000 188.840000 146.820000 189.920000 ;
      RECT 58.620000 188.840000 101.820000 189.920000 ;
      RECT 13.620000 188.840000 56.820000 189.920000 ;
      RECT 7.060000 188.840000 11.820000 189.920000 ;
      RECT 0.000000 188.840000 5.260000 189.920000 ;
      RECT 0.000000 187.200000 550.160000 188.840000 ;
      RECT 547.100000 186.200000 550.160000 187.200000 ;
      RECT 547.100000 186.120000 548.960000 186.200000 ;
      RECT 506.620000 186.120000 545.300000 187.200000 ;
      RECT 461.620000 186.120000 504.820000 187.200000 ;
      RECT 416.620000 186.120000 459.820000 187.200000 ;
      RECT 371.620000 186.120000 414.820000 187.200000 ;
      RECT 326.620000 186.120000 369.820000 187.200000 ;
      RECT 281.620000 186.120000 324.820000 187.200000 ;
      RECT 236.620000 186.120000 279.820000 187.200000 ;
      RECT 191.620000 186.120000 234.820000 187.200000 ;
      RECT 146.620000 186.120000 189.820000 187.200000 ;
      RECT 101.620000 186.120000 144.820000 187.200000 ;
      RECT 56.620000 186.120000 99.820000 187.200000 ;
      RECT 11.620000 186.120000 54.820000 187.200000 ;
      RECT 4.860000 186.120000 9.655000 187.200000 ;
      RECT 0.000000 186.120000 3.060000 187.200000 ;
      RECT 0.000000 185.220000 548.960000 186.120000 ;
      RECT 0.000000 184.480000 550.160000 185.220000 ;
      RECT 544.900000 183.400000 550.160000 184.480000 ;
      RECT 508.620000 183.400000 543.100000 184.480000 ;
      RECT 463.620000 183.400000 506.820000 184.480000 ;
      RECT 418.620000 183.400000 461.820000 184.480000 ;
      RECT 373.620000 183.400000 416.820000 184.480000 ;
      RECT 328.620000 183.400000 371.820000 184.480000 ;
      RECT 283.620000 183.400000 326.820000 184.480000 ;
      RECT 238.620000 183.400000 281.820000 184.480000 ;
      RECT 193.620000 183.400000 236.820000 184.480000 ;
      RECT 148.620000 183.400000 191.820000 184.480000 ;
      RECT 103.620000 183.400000 146.820000 184.480000 ;
      RECT 58.620000 183.400000 101.820000 184.480000 ;
      RECT 13.620000 183.400000 56.820000 184.480000 ;
      RECT 7.060000 183.400000 11.820000 184.480000 ;
      RECT 0.000000 183.400000 5.260000 184.480000 ;
      RECT 0.000000 182.540000 550.160000 183.400000 ;
      RECT 0.000000 181.760000 548.960000 182.540000 ;
      RECT 547.100000 181.560000 548.960000 181.760000 ;
      RECT 547.100000 180.680000 550.160000 181.560000 ;
      RECT 506.620000 180.680000 545.300000 181.760000 ;
      RECT 461.620000 180.680000 504.820000 181.760000 ;
      RECT 416.620000 180.680000 459.820000 181.760000 ;
      RECT 371.620000 180.680000 414.820000 181.760000 ;
      RECT 326.620000 180.680000 369.820000 181.760000 ;
      RECT 281.620000 180.680000 324.820000 181.760000 ;
      RECT 236.620000 180.680000 279.820000 181.760000 ;
      RECT 191.620000 180.680000 234.820000 181.760000 ;
      RECT 146.620000 180.680000 189.820000 181.760000 ;
      RECT 101.620000 180.680000 144.820000 181.760000 ;
      RECT 56.620000 180.680000 99.820000 181.760000 ;
      RECT 11.620000 180.680000 54.820000 181.760000 ;
      RECT 4.860000 180.680000 9.655000 181.760000 ;
      RECT 0.000000 180.680000 3.060000 181.760000 ;
      RECT 0.000000 179.490000 550.160000 180.680000 ;
      RECT 0.000000 179.040000 548.960000 179.490000 ;
      RECT 544.900000 178.510000 548.960000 179.040000 ;
      RECT 544.900000 177.960000 550.160000 178.510000 ;
      RECT 508.620000 177.960000 543.100000 179.040000 ;
      RECT 463.620000 177.960000 506.820000 179.040000 ;
      RECT 418.620000 177.960000 461.820000 179.040000 ;
      RECT 373.620000 177.960000 416.820000 179.040000 ;
      RECT 328.620000 177.960000 371.820000 179.040000 ;
      RECT 283.620000 177.960000 326.820000 179.040000 ;
      RECT 238.620000 177.960000 281.820000 179.040000 ;
      RECT 193.620000 177.960000 236.820000 179.040000 ;
      RECT 148.620000 177.960000 191.820000 179.040000 ;
      RECT 103.620000 177.960000 146.820000 179.040000 ;
      RECT 58.620000 177.960000 101.820000 179.040000 ;
      RECT 13.620000 177.960000 56.820000 179.040000 ;
      RECT 7.060000 177.960000 11.820000 179.040000 ;
      RECT 0.000000 177.960000 5.260000 179.040000 ;
      RECT 0.000000 176.320000 550.160000 177.960000 ;
      RECT 547.100000 175.830000 550.160000 176.320000 ;
      RECT 547.100000 175.240000 548.960000 175.830000 ;
      RECT 506.620000 175.240000 545.300000 176.320000 ;
      RECT 461.620000 175.240000 504.820000 176.320000 ;
      RECT 416.620000 175.240000 459.820000 176.320000 ;
      RECT 371.620000 175.240000 414.820000 176.320000 ;
      RECT 326.620000 175.240000 369.820000 176.320000 ;
      RECT 281.620000 175.240000 324.820000 176.320000 ;
      RECT 236.620000 175.240000 279.820000 176.320000 ;
      RECT 191.620000 175.240000 234.820000 176.320000 ;
      RECT 146.620000 175.240000 189.820000 176.320000 ;
      RECT 101.620000 175.240000 144.820000 176.320000 ;
      RECT 56.620000 175.240000 99.820000 176.320000 ;
      RECT 11.620000 175.240000 54.820000 176.320000 ;
      RECT 4.860000 175.240000 9.655000 176.320000 ;
      RECT 0.000000 175.240000 3.060000 176.320000 ;
      RECT 0.000000 174.850000 548.960000 175.240000 ;
      RECT 0.000000 173.600000 550.160000 174.850000 ;
      RECT 544.900000 172.520000 550.160000 173.600000 ;
      RECT 508.620000 172.520000 543.100000 173.600000 ;
      RECT 463.620000 172.520000 506.820000 173.600000 ;
      RECT 418.620000 172.520000 461.820000 173.600000 ;
      RECT 373.620000 172.520000 416.820000 173.600000 ;
      RECT 328.620000 172.520000 371.820000 173.600000 ;
      RECT 283.620000 172.520000 326.820000 173.600000 ;
      RECT 238.620000 172.520000 281.820000 173.600000 ;
      RECT 193.620000 172.520000 236.820000 173.600000 ;
      RECT 148.620000 172.520000 191.820000 173.600000 ;
      RECT 103.620000 172.520000 146.820000 173.600000 ;
      RECT 58.620000 172.520000 101.820000 173.600000 ;
      RECT 13.620000 172.520000 56.820000 173.600000 ;
      RECT 7.060000 172.520000 11.820000 173.600000 ;
      RECT 0.000000 172.520000 5.260000 173.600000 ;
      RECT 0.000000 172.170000 550.160000 172.520000 ;
      RECT 0.000000 171.190000 548.960000 172.170000 ;
      RECT 0.000000 170.880000 550.160000 171.190000 ;
      RECT 547.100000 169.800000 550.160000 170.880000 ;
      RECT 506.620000 169.800000 545.300000 170.880000 ;
      RECT 461.620000 169.800000 504.820000 170.880000 ;
      RECT 416.620000 169.800000 459.820000 170.880000 ;
      RECT 371.620000 169.800000 414.820000 170.880000 ;
      RECT 326.620000 169.800000 369.820000 170.880000 ;
      RECT 281.620000 169.800000 324.820000 170.880000 ;
      RECT 236.620000 169.800000 279.820000 170.880000 ;
      RECT 191.620000 169.800000 234.820000 170.880000 ;
      RECT 146.620000 169.800000 189.820000 170.880000 ;
      RECT 101.620000 169.800000 144.820000 170.880000 ;
      RECT 56.620000 169.800000 99.820000 170.880000 ;
      RECT 11.620000 169.800000 54.820000 170.880000 ;
      RECT 4.860000 169.800000 9.655000 170.880000 ;
      RECT 0.000000 169.800000 3.060000 170.880000 ;
      RECT 0.000000 169.120000 550.160000 169.800000 ;
      RECT 0.000000 168.160000 548.960000 169.120000 ;
      RECT 544.900000 168.140000 548.960000 168.160000 ;
      RECT 544.900000 167.080000 550.160000 168.140000 ;
      RECT 508.620000 167.080000 543.100000 168.160000 ;
      RECT 463.620000 167.080000 506.820000 168.160000 ;
      RECT 418.620000 167.080000 461.820000 168.160000 ;
      RECT 373.620000 167.080000 416.820000 168.160000 ;
      RECT 328.620000 167.080000 371.820000 168.160000 ;
      RECT 283.620000 167.080000 326.820000 168.160000 ;
      RECT 238.620000 167.080000 281.820000 168.160000 ;
      RECT 193.620000 167.080000 236.820000 168.160000 ;
      RECT 148.620000 167.080000 191.820000 168.160000 ;
      RECT 103.620000 167.080000 146.820000 168.160000 ;
      RECT 58.620000 167.080000 101.820000 168.160000 ;
      RECT 13.620000 167.080000 56.820000 168.160000 ;
      RECT 7.060000 167.080000 11.820000 168.160000 ;
      RECT 0.000000 167.080000 5.260000 168.160000 ;
      RECT 0.000000 165.460000 550.160000 167.080000 ;
      RECT 0.000000 165.440000 548.960000 165.460000 ;
      RECT 547.100000 164.480000 548.960000 165.440000 ;
      RECT 547.100000 164.360000 550.160000 164.480000 ;
      RECT 506.620000 164.360000 545.300000 165.440000 ;
      RECT 461.620000 164.360000 504.820000 165.440000 ;
      RECT 416.620000 164.360000 459.820000 165.440000 ;
      RECT 371.620000 164.360000 414.820000 165.440000 ;
      RECT 326.620000 164.360000 369.820000 165.440000 ;
      RECT 281.620000 164.360000 324.820000 165.440000 ;
      RECT 236.620000 164.360000 279.820000 165.440000 ;
      RECT 191.620000 164.360000 234.820000 165.440000 ;
      RECT 146.620000 164.360000 189.820000 165.440000 ;
      RECT 101.620000 164.360000 144.820000 165.440000 ;
      RECT 56.620000 164.360000 99.820000 165.440000 ;
      RECT 11.620000 164.360000 54.820000 165.440000 ;
      RECT 4.860000 164.360000 9.655000 165.440000 ;
      RECT 0.000000 164.360000 3.060000 165.440000 ;
      RECT 0.000000 162.720000 550.160000 164.360000 ;
      RECT 544.900000 161.800000 550.160000 162.720000 ;
      RECT 544.900000 161.640000 548.960000 161.800000 ;
      RECT 508.620000 161.640000 543.100000 162.720000 ;
      RECT 463.620000 161.640000 506.820000 162.720000 ;
      RECT 418.620000 161.640000 461.820000 162.720000 ;
      RECT 373.620000 161.640000 416.820000 162.720000 ;
      RECT 328.620000 161.640000 371.820000 162.720000 ;
      RECT 283.620000 161.640000 326.820000 162.720000 ;
      RECT 238.620000 161.640000 281.820000 162.720000 ;
      RECT 193.620000 161.640000 236.820000 162.720000 ;
      RECT 148.620000 161.640000 191.820000 162.720000 ;
      RECT 103.620000 161.640000 146.820000 162.720000 ;
      RECT 58.620000 161.640000 101.820000 162.720000 ;
      RECT 13.620000 161.640000 56.820000 162.720000 ;
      RECT 7.060000 161.640000 11.820000 162.720000 ;
      RECT 0.000000 161.640000 5.260000 162.720000 ;
      RECT 0.000000 160.820000 548.960000 161.640000 ;
      RECT 0.000000 160.000000 550.160000 160.820000 ;
      RECT 547.100000 158.920000 550.160000 160.000000 ;
      RECT 506.620000 158.920000 545.300000 160.000000 ;
      RECT 461.620000 158.920000 504.820000 160.000000 ;
      RECT 416.620000 158.920000 459.820000 160.000000 ;
      RECT 371.620000 158.920000 414.820000 160.000000 ;
      RECT 326.620000 158.920000 369.820000 160.000000 ;
      RECT 281.620000 158.920000 324.820000 160.000000 ;
      RECT 236.620000 158.920000 279.820000 160.000000 ;
      RECT 191.620000 158.920000 234.820000 160.000000 ;
      RECT 146.620000 158.920000 189.820000 160.000000 ;
      RECT 101.620000 158.920000 144.820000 160.000000 ;
      RECT 56.620000 158.920000 99.820000 160.000000 ;
      RECT 11.620000 158.920000 54.820000 160.000000 ;
      RECT 4.860000 158.920000 9.655000 160.000000 ;
      RECT 0.000000 158.920000 3.060000 160.000000 ;
      RECT 0.000000 158.750000 550.160000 158.920000 ;
      RECT 0.000000 157.770000 548.960000 158.750000 ;
      RECT 0.000000 157.280000 550.160000 157.770000 ;
      RECT 544.900000 156.200000 550.160000 157.280000 ;
      RECT 508.620000 156.200000 543.100000 157.280000 ;
      RECT 463.620000 156.200000 506.820000 157.280000 ;
      RECT 418.620000 156.200000 461.820000 157.280000 ;
      RECT 373.620000 156.200000 416.820000 157.280000 ;
      RECT 328.620000 156.200000 371.820000 157.280000 ;
      RECT 283.620000 156.200000 326.820000 157.280000 ;
      RECT 238.620000 156.200000 281.820000 157.280000 ;
      RECT 193.620000 156.200000 236.820000 157.280000 ;
      RECT 148.620000 156.200000 191.820000 157.280000 ;
      RECT 103.620000 156.200000 146.820000 157.280000 ;
      RECT 58.620000 156.200000 101.820000 157.280000 ;
      RECT 13.620000 156.200000 56.820000 157.280000 ;
      RECT 7.060000 156.200000 11.820000 157.280000 ;
      RECT 0.000000 156.200000 5.260000 157.280000 ;
      RECT 0.000000 155.090000 550.160000 156.200000 ;
      RECT 0.000000 154.560000 548.960000 155.090000 ;
      RECT 547.100000 154.110000 548.960000 154.560000 ;
      RECT 547.100000 153.480000 550.160000 154.110000 ;
      RECT 506.620000 153.480000 545.300000 154.560000 ;
      RECT 461.620000 153.480000 504.820000 154.560000 ;
      RECT 416.620000 153.480000 459.820000 154.560000 ;
      RECT 371.620000 153.480000 414.820000 154.560000 ;
      RECT 326.620000 153.480000 369.820000 154.560000 ;
      RECT 281.620000 153.480000 324.820000 154.560000 ;
      RECT 236.620000 153.480000 279.820000 154.560000 ;
      RECT 191.620000 153.480000 234.820000 154.560000 ;
      RECT 146.620000 153.480000 189.820000 154.560000 ;
      RECT 101.620000 153.480000 144.820000 154.560000 ;
      RECT 56.620000 153.480000 99.820000 154.560000 ;
      RECT 11.620000 153.480000 54.820000 154.560000 ;
      RECT 4.860000 153.480000 9.655000 154.560000 ;
      RECT 0.000000 153.480000 3.060000 154.560000 ;
      RECT 0.000000 151.840000 550.160000 153.480000 ;
      RECT 544.900000 151.430000 550.160000 151.840000 ;
      RECT 544.900000 150.760000 548.960000 151.430000 ;
      RECT 508.620000 150.760000 543.100000 151.840000 ;
      RECT 463.620000 150.760000 506.820000 151.840000 ;
      RECT 418.620000 150.760000 461.820000 151.840000 ;
      RECT 373.620000 150.760000 416.820000 151.840000 ;
      RECT 328.620000 150.760000 371.820000 151.840000 ;
      RECT 283.620000 150.760000 326.820000 151.840000 ;
      RECT 238.620000 150.760000 281.820000 151.840000 ;
      RECT 193.620000 150.760000 236.820000 151.840000 ;
      RECT 148.620000 150.760000 191.820000 151.840000 ;
      RECT 103.620000 150.760000 146.820000 151.840000 ;
      RECT 58.620000 150.760000 101.820000 151.840000 ;
      RECT 13.620000 150.760000 56.820000 151.840000 ;
      RECT 7.060000 150.760000 11.820000 151.840000 ;
      RECT 0.000000 150.760000 5.260000 151.840000 ;
      RECT 0.000000 150.450000 548.960000 150.760000 ;
      RECT 0.000000 149.120000 550.160000 150.450000 ;
      RECT 547.100000 148.380000 550.160000 149.120000 ;
      RECT 547.100000 148.040000 548.960000 148.380000 ;
      RECT 506.620000 148.040000 545.300000 149.120000 ;
      RECT 461.620000 148.040000 504.820000 149.120000 ;
      RECT 416.620000 148.040000 459.820000 149.120000 ;
      RECT 371.620000 148.040000 414.820000 149.120000 ;
      RECT 326.620000 148.040000 369.820000 149.120000 ;
      RECT 281.620000 148.040000 324.820000 149.120000 ;
      RECT 236.620000 148.040000 279.820000 149.120000 ;
      RECT 191.620000 148.040000 234.820000 149.120000 ;
      RECT 146.620000 148.040000 189.820000 149.120000 ;
      RECT 101.620000 148.040000 144.820000 149.120000 ;
      RECT 56.620000 148.040000 99.820000 149.120000 ;
      RECT 11.620000 148.040000 54.820000 149.120000 ;
      RECT 4.860000 148.040000 9.655000 149.120000 ;
      RECT 0.000000 148.040000 3.060000 149.120000 ;
      RECT 0.000000 147.400000 548.960000 148.040000 ;
      RECT 0.000000 146.400000 550.160000 147.400000 ;
      RECT 544.900000 145.320000 550.160000 146.400000 ;
      RECT 508.620000 145.320000 543.100000 146.400000 ;
      RECT 463.620000 145.320000 506.820000 146.400000 ;
      RECT 418.620000 145.320000 461.820000 146.400000 ;
      RECT 373.620000 145.320000 416.820000 146.400000 ;
      RECT 328.620000 145.320000 371.820000 146.400000 ;
      RECT 283.620000 145.320000 326.820000 146.400000 ;
      RECT 238.620000 145.320000 281.820000 146.400000 ;
      RECT 193.620000 145.320000 236.820000 146.400000 ;
      RECT 148.620000 145.320000 191.820000 146.400000 ;
      RECT 103.620000 145.320000 146.820000 146.400000 ;
      RECT 58.620000 145.320000 101.820000 146.400000 ;
      RECT 13.620000 145.320000 56.820000 146.400000 ;
      RECT 7.060000 145.320000 11.820000 146.400000 ;
      RECT 0.000000 145.320000 5.260000 146.400000 ;
      RECT 0.000000 144.720000 550.160000 145.320000 ;
      RECT 0.000000 143.740000 548.960000 144.720000 ;
      RECT 0.000000 143.680000 550.160000 143.740000 ;
      RECT 547.100000 142.600000 550.160000 143.680000 ;
      RECT 506.620000 142.600000 545.300000 143.680000 ;
      RECT 461.620000 142.600000 504.820000 143.680000 ;
      RECT 416.620000 142.600000 459.820000 143.680000 ;
      RECT 371.620000 142.600000 414.820000 143.680000 ;
      RECT 326.620000 142.600000 369.820000 143.680000 ;
      RECT 281.620000 142.600000 324.820000 143.680000 ;
      RECT 236.620000 142.600000 279.820000 143.680000 ;
      RECT 191.620000 142.600000 234.820000 143.680000 ;
      RECT 146.620000 142.600000 189.820000 143.680000 ;
      RECT 101.620000 142.600000 144.820000 143.680000 ;
      RECT 56.620000 142.600000 99.820000 143.680000 ;
      RECT 11.620000 142.600000 54.820000 143.680000 ;
      RECT 4.860000 142.600000 9.655000 143.680000 ;
      RECT 0.000000 142.600000 3.060000 143.680000 ;
      RECT 0.000000 141.060000 550.160000 142.600000 ;
      RECT 0.000000 140.960000 548.960000 141.060000 ;
      RECT 544.900000 140.080000 548.960000 140.960000 ;
      RECT 544.900000 139.880000 550.160000 140.080000 ;
      RECT 508.620000 139.880000 543.100000 140.960000 ;
      RECT 463.620000 139.880000 506.820000 140.960000 ;
      RECT 418.620000 139.880000 461.820000 140.960000 ;
      RECT 373.620000 139.880000 416.820000 140.960000 ;
      RECT 328.620000 139.880000 371.820000 140.960000 ;
      RECT 283.620000 139.880000 326.820000 140.960000 ;
      RECT 238.620000 139.880000 281.820000 140.960000 ;
      RECT 193.620000 139.880000 236.820000 140.960000 ;
      RECT 148.620000 139.880000 191.820000 140.960000 ;
      RECT 103.620000 139.880000 146.820000 140.960000 ;
      RECT 58.620000 139.880000 101.820000 140.960000 ;
      RECT 13.620000 139.880000 56.820000 140.960000 ;
      RECT 7.060000 139.880000 11.820000 140.960000 ;
      RECT 0.000000 139.880000 5.260000 140.960000 ;
      RECT 0.000000 138.240000 550.160000 139.880000 ;
      RECT 547.100000 138.010000 550.160000 138.240000 ;
      RECT 547.100000 137.160000 548.960000 138.010000 ;
      RECT 506.620000 137.160000 545.300000 138.240000 ;
      RECT 461.620000 137.160000 504.820000 138.240000 ;
      RECT 416.620000 137.160000 459.820000 138.240000 ;
      RECT 371.620000 137.160000 414.820000 138.240000 ;
      RECT 326.620000 137.160000 369.820000 138.240000 ;
      RECT 281.620000 137.160000 324.820000 138.240000 ;
      RECT 236.620000 137.160000 279.820000 138.240000 ;
      RECT 191.620000 137.160000 234.820000 138.240000 ;
      RECT 146.620000 137.160000 189.820000 138.240000 ;
      RECT 101.620000 137.160000 144.820000 138.240000 ;
      RECT 56.620000 137.160000 99.820000 138.240000 ;
      RECT 11.620000 137.160000 54.820000 138.240000 ;
      RECT 4.860000 137.160000 9.655000 138.240000 ;
      RECT 0.000000 137.160000 3.060000 138.240000 ;
      RECT 0.000000 137.030000 548.960000 137.160000 ;
      RECT 0.000000 135.520000 550.160000 137.030000 ;
      RECT 544.900000 134.440000 550.160000 135.520000 ;
      RECT 508.620000 134.440000 543.100000 135.520000 ;
      RECT 463.620000 134.440000 506.820000 135.520000 ;
      RECT 418.620000 134.440000 461.820000 135.520000 ;
      RECT 373.620000 134.440000 416.820000 135.520000 ;
      RECT 328.620000 134.440000 371.820000 135.520000 ;
      RECT 283.620000 134.440000 326.820000 135.520000 ;
      RECT 238.620000 134.440000 281.820000 135.520000 ;
      RECT 193.620000 134.440000 236.820000 135.520000 ;
      RECT 148.620000 134.440000 191.820000 135.520000 ;
      RECT 103.620000 134.440000 146.820000 135.520000 ;
      RECT 58.620000 134.440000 101.820000 135.520000 ;
      RECT 13.620000 134.440000 56.820000 135.520000 ;
      RECT 7.060000 134.440000 11.820000 135.520000 ;
      RECT 0.000000 134.440000 5.260000 135.520000 ;
      RECT 0.000000 134.350000 550.160000 134.440000 ;
      RECT 0.000000 133.370000 548.960000 134.350000 ;
      RECT 0.000000 132.800000 550.160000 133.370000 ;
      RECT 547.100000 131.720000 550.160000 132.800000 ;
      RECT 506.620000 131.720000 545.300000 132.800000 ;
      RECT 461.620000 131.720000 504.820000 132.800000 ;
      RECT 416.620000 131.720000 459.820000 132.800000 ;
      RECT 371.620000 131.720000 414.820000 132.800000 ;
      RECT 326.620000 131.720000 369.820000 132.800000 ;
      RECT 281.620000 131.720000 324.820000 132.800000 ;
      RECT 236.620000 131.720000 279.820000 132.800000 ;
      RECT 191.620000 131.720000 234.820000 132.800000 ;
      RECT 146.620000 131.720000 189.820000 132.800000 ;
      RECT 101.620000 131.720000 144.820000 132.800000 ;
      RECT 56.620000 131.720000 99.820000 132.800000 ;
      RECT 11.620000 131.720000 54.820000 132.800000 ;
      RECT 4.860000 131.720000 9.655000 132.800000 ;
      RECT 0.000000 131.720000 3.060000 132.800000 ;
      RECT 0.000000 130.690000 550.160000 131.720000 ;
      RECT 0.000000 130.080000 548.960000 130.690000 ;
      RECT 544.900000 129.710000 548.960000 130.080000 ;
      RECT 544.900000 129.000000 550.160000 129.710000 ;
      RECT 508.620000 129.000000 543.100000 130.080000 ;
      RECT 463.620000 129.000000 506.820000 130.080000 ;
      RECT 418.620000 129.000000 461.820000 130.080000 ;
      RECT 373.620000 129.000000 416.820000 130.080000 ;
      RECT 328.620000 129.000000 371.820000 130.080000 ;
      RECT 283.620000 129.000000 326.820000 130.080000 ;
      RECT 238.620000 129.000000 281.820000 130.080000 ;
      RECT 193.620000 129.000000 236.820000 130.080000 ;
      RECT 148.620000 129.000000 191.820000 130.080000 ;
      RECT 103.620000 129.000000 146.820000 130.080000 ;
      RECT 58.620000 129.000000 101.820000 130.080000 ;
      RECT 13.620000 129.000000 56.820000 130.080000 ;
      RECT 7.060000 129.000000 11.820000 130.080000 ;
      RECT 0.000000 129.000000 5.260000 130.080000 ;
      RECT 0.000000 127.640000 550.160000 129.000000 ;
      RECT 0.000000 127.360000 548.960000 127.640000 ;
      RECT 547.100000 126.660000 548.960000 127.360000 ;
      RECT 547.100000 126.280000 550.160000 126.660000 ;
      RECT 506.620000 126.280000 545.300000 127.360000 ;
      RECT 461.620000 126.280000 504.820000 127.360000 ;
      RECT 416.620000 126.280000 459.820000 127.360000 ;
      RECT 371.620000 126.280000 414.820000 127.360000 ;
      RECT 326.620000 126.280000 369.820000 127.360000 ;
      RECT 281.620000 126.280000 324.820000 127.360000 ;
      RECT 236.620000 126.280000 279.820000 127.360000 ;
      RECT 191.620000 126.280000 234.820000 127.360000 ;
      RECT 146.620000 126.280000 189.820000 127.360000 ;
      RECT 101.620000 126.280000 144.820000 127.360000 ;
      RECT 56.620000 126.280000 99.820000 127.360000 ;
      RECT 11.620000 126.280000 54.820000 127.360000 ;
      RECT 4.860000 126.280000 9.655000 127.360000 ;
      RECT 0.000000 126.280000 3.060000 127.360000 ;
      RECT 0.000000 124.640000 550.160000 126.280000 ;
      RECT 544.900000 123.980000 550.160000 124.640000 ;
      RECT 544.900000 123.560000 548.960000 123.980000 ;
      RECT 508.620000 123.560000 543.100000 124.640000 ;
      RECT 463.620000 123.560000 506.820000 124.640000 ;
      RECT 418.620000 123.560000 461.820000 124.640000 ;
      RECT 373.620000 123.560000 416.820000 124.640000 ;
      RECT 328.620000 123.560000 371.820000 124.640000 ;
      RECT 283.620000 123.560000 326.820000 124.640000 ;
      RECT 238.620000 123.560000 281.820000 124.640000 ;
      RECT 193.620000 123.560000 236.820000 124.640000 ;
      RECT 148.620000 123.560000 191.820000 124.640000 ;
      RECT 103.620000 123.560000 146.820000 124.640000 ;
      RECT 58.620000 123.560000 101.820000 124.640000 ;
      RECT 13.620000 123.560000 56.820000 124.640000 ;
      RECT 7.060000 123.560000 11.820000 124.640000 ;
      RECT 0.000000 123.560000 5.260000 124.640000 ;
      RECT 0.000000 123.000000 548.960000 123.560000 ;
      RECT 0.000000 121.920000 550.160000 123.000000 ;
      RECT 547.100000 120.840000 550.160000 121.920000 ;
      RECT 506.620000 120.840000 545.300000 121.920000 ;
      RECT 461.620000 120.840000 504.820000 121.920000 ;
      RECT 416.620000 120.840000 459.820000 121.920000 ;
      RECT 371.620000 120.840000 414.820000 121.920000 ;
      RECT 326.620000 120.840000 369.820000 121.920000 ;
      RECT 281.620000 120.840000 324.820000 121.920000 ;
      RECT 236.620000 120.840000 279.820000 121.920000 ;
      RECT 191.620000 120.840000 234.820000 121.920000 ;
      RECT 146.620000 120.840000 189.820000 121.920000 ;
      RECT 101.620000 120.840000 144.820000 121.920000 ;
      RECT 56.620000 120.840000 99.820000 121.920000 ;
      RECT 11.620000 120.840000 54.820000 121.920000 ;
      RECT 4.860000 120.840000 9.655000 121.920000 ;
      RECT 0.000000 120.840000 3.060000 121.920000 ;
      RECT 0.000000 120.320000 550.160000 120.840000 ;
      RECT 0.000000 119.340000 548.960000 120.320000 ;
      RECT 0.000000 119.200000 550.160000 119.340000 ;
      RECT 544.900000 118.120000 550.160000 119.200000 ;
      RECT 508.620000 118.120000 543.100000 119.200000 ;
      RECT 463.620000 118.120000 506.820000 119.200000 ;
      RECT 418.620000 118.120000 461.820000 119.200000 ;
      RECT 373.620000 118.120000 416.820000 119.200000 ;
      RECT 328.620000 118.120000 371.820000 119.200000 ;
      RECT 283.620000 118.120000 326.820000 119.200000 ;
      RECT 238.620000 118.120000 281.820000 119.200000 ;
      RECT 193.620000 118.120000 236.820000 119.200000 ;
      RECT 148.620000 118.120000 191.820000 119.200000 ;
      RECT 103.620000 118.120000 146.820000 119.200000 ;
      RECT 58.620000 118.120000 101.820000 119.200000 ;
      RECT 13.620000 118.120000 56.820000 119.200000 ;
      RECT 7.060000 118.120000 11.820000 119.200000 ;
      RECT 0.000000 118.120000 5.260000 119.200000 ;
      RECT 0.000000 117.270000 550.160000 118.120000 ;
      RECT 0.000000 116.480000 548.960000 117.270000 ;
      RECT 547.100000 116.290000 548.960000 116.480000 ;
      RECT 547.100000 115.400000 550.160000 116.290000 ;
      RECT 506.620000 115.400000 545.300000 116.480000 ;
      RECT 461.620000 115.400000 504.820000 116.480000 ;
      RECT 416.620000 115.400000 459.820000 116.480000 ;
      RECT 371.620000 115.400000 414.820000 116.480000 ;
      RECT 326.620000 115.400000 369.820000 116.480000 ;
      RECT 281.620000 115.400000 324.820000 116.480000 ;
      RECT 236.620000 115.400000 279.820000 116.480000 ;
      RECT 191.620000 115.400000 234.820000 116.480000 ;
      RECT 146.620000 115.400000 189.820000 116.480000 ;
      RECT 101.620000 115.400000 144.820000 116.480000 ;
      RECT 56.620000 115.400000 99.820000 116.480000 ;
      RECT 11.620000 115.400000 54.820000 116.480000 ;
      RECT 4.860000 115.400000 9.655000 116.480000 ;
      RECT 0.000000 115.400000 3.060000 116.480000 ;
      RECT 0.000000 113.760000 550.160000 115.400000 ;
      RECT 544.900000 113.610000 550.160000 113.760000 ;
      RECT 544.900000 112.680000 548.960000 113.610000 ;
      RECT 508.620000 112.680000 543.100000 113.760000 ;
      RECT 463.620000 112.680000 506.820000 113.760000 ;
      RECT 418.620000 112.680000 461.820000 113.760000 ;
      RECT 373.620000 112.680000 416.820000 113.760000 ;
      RECT 328.620000 112.680000 371.820000 113.760000 ;
      RECT 283.620000 112.680000 326.820000 113.760000 ;
      RECT 238.620000 112.680000 281.820000 113.760000 ;
      RECT 193.620000 112.680000 236.820000 113.760000 ;
      RECT 148.620000 112.680000 191.820000 113.760000 ;
      RECT 103.620000 112.680000 146.820000 113.760000 ;
      RECT 58.620000 112.680000 101.820000 113.760000 ;
      RECT 13.620000 112.680000 56.820000 113.760000 ;
      RECT 7.060000 112.680000 11.820000 113.760000 ;
      RECT 0.000000 112.680000 5.260000 113.760000 ;
      RECT 0.000000 112.630000 548.960000 112.680000 ;
      RECT 0.000000 111.040000 550.160000 112.630000 ;
      RECT 547.100000 109.960000 550.160000 111.040000 ;
      RECT 506.620000 109.960000 545.300000 111.040000 ;
      RECT 461.620000 109.960000 504.820000 111.040000 ;
      RECT 416.620000 109.960000 459.820000 111.040000 ;
      RECT 371.620000 109.960000 414.820000 111.040000 ;
      RECT 326.620000 109.960000 369.820000 111.040000 ;
      RECT 281.620000 109.960000 324.820000 111.040000 ;
      RECT 236.620000 109.960000 279.820000 111.040000 ;
      RECT 191.620000 109.960000 234.820000 111.040000 ;
      RECT 146.620000 109.960000 189.820000 111.040000 ;
      RECT 101.620000 109.960000 144.820000 111.040000 ;
      RECT 56.620000 109.960000 99.820000 111.040000 ;
      RECT 11.620000 109.960000 54.820000 111.040000 ;
      RECT 4.860000 109.960000 9.655000 111.040000 ;
      RECT 0.000000 109.960000 3.060000 111.040000 ;
      RECT 0.000000 109.950000 550.160000 109.960000 ;
      RECT 0.000000 108.970000 548.960000 109.950000 ;
      RECT 0.000000 108.320000 550.160000 108.970000 ;
      RECT 544.900000 107.240000 550.160000 108.320000 ;
      RECT 508.620000 107.240000 543.100000 108.320000 ;
      RECT 463.620000 107.240000 506.820000 108.320000 ;
      RECT 418.620000 107.240000 461.820000 108.320000 ;
      RECT 373.620000 107.240000 416.820000 108.320000 ;
      RECT 328.620000 107.240000 371.820000 108.320000 ;
      RECT 283.620000 107.240000 326.820000 108.320000 ;
      RECT 238.620000 107.240000 281.820000 108.320000 ;
      RECT 193.620000 107.240000 236.820000 108.320000 ;
      RECT 148.620000 107.240000 191.820000 108.320000 ;
      RECT 103.620000 107.240000 146.820000 108.320000 ;
      RECT 58.620000 107.240000 101.820000 108.320000 ;
      RECT 13.620000 107.240000 56.820000 108.320000 ;
      RECT 7.060000 107.240000 11.820000 108.320000 ;
      RECT 0.000000 107.240000 5.260000 108.320000 ;
      RECT 0.000000 106.900000 550.160000 107.240000 ;
      RECT 0.000000 105.920000 548.960000 106.900000 ;
      RECT 0.000000 105.600000 550.160000 105.920000 ;
      RECT 547.100000 104.520000 550.160000 105.600000 ;
      RECT 506.620000 104.520000 545.300000 105.600000 ;
      RECT 461.620000 104.520000 504.820000 105.600000 ;
      RECT 416.620000 104.520000 459.820000 105.600000 ;
      RECT 371.620000 104.520000 414.820000 105.600000 ;
      RECT 326.620000 104.520000 369.820000 105.600000 ;
      RECT 281.620000 104.520000 324.820000 105.600000 ;
      RECT 236.620000 104.520000 279.820000 105.600000 ;
      RECT 191.620000 104.520000 234.820000 105.600000 ;
      RECT 146.620000 104.520000 189.820000 105.600000 ;
      RECT 101.620000 104.520000 144.820000 105.600000 ;
      RECT 56.620000 104.520000 99.820000 105.600000 ;
      RECT 11.620000 104.520000 54.820000 105.600000 ;
      RECT 4.860000 104.520000 9.655000 105.600000 ;
      RECT 0.000000 104.520000 3.060000 105.600000 ;
      RECT 0.000000 103.240000 550.160000 104.520000 ;
      RECT 0.000000 102.880000 548.960000 103.240000 ;
      RECT 544.900000 102.260000 548.960000 102.880000 ;
      RECT 544.900000 101.800000 550.160000 102.260000 ;
      RECT 508.620000 101.800000 543.100000 102.880000 ;
      RECT 463.620000 101.800000 506.820000 102.880000 ;
      RECT 418.620000 101.800000 461.820000 102.880000 ;
      RECT 373.620000 101.800000 416.820000 102.880000 ;
      RECT 328.620000 101.800000 371.820000 102.880000 ;
      RECT 283.620000 101.800000 326.820000 102.880000 ;
      RECT 238.620000 101.800000 281.820000 102.880000 ;
      RECT 193.620000 101.800000 236.820000 102.880000 ;
      RECT 148.620000 101.800000 191.820000 102.880000 ;
      RECT 103.620000 101.800000 146.820000 102.880000 ;
      RECT 58.620000 101.800000 101.820000 102.880000 ;
      RECT 13.620000 101.800000 56.820000 102.880000 ;
      RECT 7.060000 101.800000 11.820000 102.880000 ;
      RECT 0.000000 101.800000 5.260000 102.880000 ;
      RECT 0.000000 100.190000 550.160000 101.800000 ;
      RECT 0.000000 100.160000 548.960000 100.190000 ;
      RECT 547.100000 99.210000 548.960000 100.160000 ;
      RECT 547.100000 99.080000 550.160000 99.210000 ;
      RECT 506.620000 99.080000 545.300000 100.160000 ;
      RECT 461.620000 99.080000 504.820000 100.160000 ;
      RECT 416.620000 99.080000 459.820000 100.160000 ;
      RECT 371.620000 99.080000 414.820000 100.160000 ;
      RECT 326.620000 99.080000 369.820000 100.160000 ;
      RECT 281.620000 99.080000 324.820000 100.160000 ;
      RECT 236.620000 99.080000 279.820000 100.160000 ;
      RECT 191.620000 99.080000 234.820000 100.160000 ;
      RECT 146.620000 99.080000 189.820000 100.160000 ;
      RECT 101.620000 99.080000 144.820000 100.160000 ;
      RECT 56.620000 99.080000 99.820000 100.160000 ;
      RECT 11.620000 99.080000 54.820000 100.160000 ;
      RECT 4.860000 99.080000 9.655000 100.160000 ;
      RECT 0.000000 99.080000 3.060000 100.160000 ;
      RECT 0.000000 97.440000 550.160000 99.080000 ;
      RECT 544.900000 96.530000 550.160000 97.440000 ;
      RECT 544.900000 96.360000 548.960000 96.530000 ;
      RECT 508.620000 96.360000 543.100000 97.440000 ;
      RECT 463.620000 96.360000 506.820000 97.440000 ;
      RECT 418.620000 96.360000 461.820000 97.440000 ;
      RECT 373.620000 96.360000 416.820000 97.440000 ;
      RECT 328.620000 96.360000 371.820000 97.440000 ;
      RECT 283.620000 96.360000 326.820000 97.440000 ;
      RECT 238.620000 96.360000 281.820000 97.440000 ;
      RECT 193.620000 96.360000 236.820000 97.440000 ;
      RECT 148.620000 96.360000 191.820000 97.440000 ;
      RECT 103.620000 96.360000 146.820000 97.440000 ;
      RECT 58.620000 96.360000 101.820000 97.440000 ;
      RECT 13.620000 96.360000 56.820000 97.440000 ;
      RECT 7.060000 96.360000 11.820000 97.440000 ;
      RECT 0.000000 96.360000 5.260000 97.440000 ;
      RECT 0.000000 95.550000 548.960000 96.360000 ;
      RECT 0.000000 94.720000 550.160000 95.550000 ;
      RECT 547.100000 93.640000 550.160000 94.720000 ;
      RECT 506.620000 93.640000 545.300000 94.720000 ;
      RECT 461.620000 93.640000 504.820000 94.720000 ;
      RECT 416.620000 93.640000 459.820000 94.720000 ;
      RECT 371.620000 93.640000 414.820000 94.720000 ;
      RECT 326.620000 93.640000 369.820000 94.720000 ;
      RECT 281.620000 93.640000 324.820000 94.720000 ;
      RECT 236.620000 93.640000 279.820000 94.720000 ;
      RECT 191.620000 93.640000 234.820000 94.720000 ;
      RECT 146.620000 93.640000 189.820000 94.720000 ;
      RECT 101.620000 93.640000 144.820000 94.720000 ;
      RECT 56.620000 93.640000 99.820000 94.720000 ;
      RECT 11.620000 93.640000 54.820000 94.720000 ;
      RECT 4.860000 93.640000 9.655000 94.720000 ;
      RECT 0.000000 93.640000 3.060000 94.720000 ;
      RECT 0.000000 92.870000 550.160000 93.640000 ;
      RECT 0.000000 92.000000 548.960000 92.870000 ;
      RECT 544.900000 91.890000 548.960000 92.000000 ;
      RECT 544.900000 90.920000 550.160000 91.890000 ;
      RECT 508.620000 90.920000 543.100000 92.000000 ;
      RECT 463.620000 90.920000 506.820000 92.000000 ;
      RECT 418.620000 90.920000 461.820000 92.000000 ;
      RECT 373.620000 90.920000 416.820000 92.000000 ;
      RECT 328.620000 90.920000 371.820000 92.000000 ;
      RECT 283.620000 90.920000 326.820000 92.000000 ;
      RECT 238.620000 90.920000 281.820000 92.000000 ;
      RECT 193.620000 90.920000 236.820000 92.000000 ;
      RECT 148.620000 90.920000 191.820000 92.000000 ;
      RECT 103.620000 90.920000 146.820000 92.000000 ;
      RECT 58.620000 90.920000 101.820000 92.000000 ;
      RECT 13.620000 90.920000 56.820000 92.000000 ;
      RECT 7.060000 90.920000 11.820000 92.000000 ;
      RECT 0.000000 90.920000 5.260000 92.000000 ;
      RECT 0.000000 89.820000 550.160000 90.920000 ;
      RECT 0.000000 89.280000 548.960000 89.820000 ;
      RECT 547.100000 88.840000 548.960000 89.280000 ;
      RECT 547.100000 88.200000 550.160000 88.840000 ;
      RECT 506.620000 88.200000 545.300000 89.280000 ;
      RECT 461.620000 88.200000 504.820000 89.280000 ;
      RECT 416.620000 88.200000 459.820000 89.280000 ;
      RECT 371.620000 88.200000 414.820000 89.280000 ;
      RECT 326.620000 88.200000 369.820000 89.280000 ;
      RECT 281.620000 88.200000 324.820000 89.280000 ;
      RECT 236.620000 88.200000 279.820000 89.280000 ;
      RECT 191.620000 88.200000 234.820000 89.280000 ;
      RECT 146.620000 88.200000 189.820000 89.280000 ;
      RECT 101.620000 88.200000 144.820000 89.280000 ;
      RECT 56.620000 88.200000 99.820000 89.280000 ;
      RECT 11.620000 88.200000 54.820000 89.280000 ;
      RECT 4.860000 88.200000 9.655000 89.280000 ;
      RECT 0.000000 88.200000 3.060000 89.280000 ;
      RECT 0.000000 86.560000 550.160000 88.200000 ;
      RECT 544.900000 86.160000 550.160000 86.560000 ;
      RECT 544.900000 85.480000 548.960000 86.160000 ;
      RECT 508.620000 85.480000 543.100000 86.560000 ;
      RECT 463.620000 85.480000 506.820000 86.560000 ;
      RECT 418.620000 85.480000 461.820000 86.560000 ;
      RECT 373.620000 85.480000 416.820000 86.560000 ;
      RECT 328.620000 85.480000 371.820000 86.560000 ;
      RECT 283.620000 85.480000 326.820000 86.560000 ;
      RECT 238.620000 85.480000 281.820000 86.560000 ;
      RECT 193.620000 85.480000 236.820000 86.560000 ;
      RECT 148.620000 85.480000 191.820000 86.560000 ;
      RECT 103.620000 85.480000 146.820000 86.560000 ;
      RECT 58.620000 85.480000 101.820000 86.560000 ;
      RECT 13.620000 85.480000 56.820000 86.560000 ;
      RECT 7.060000 85.480000 11.820000 86.560000 ;
      RECT 0.000000 85.480000 5.260000 86.560000 ;
      RECT 0.000000 85.180000 548.960000 85.480000 ;
      RECT 0.000000 83.840000 550.160000 85.180000 ;
      RECT 547.100000 82.760000 550.160000 83.840000 ;
      RECT 506.620000 82.760000 545.300000 83.840000 ;
      RECT 461.620000 82.760000 504.820000 83.840000 ;
      RECT 416.620000 82.760000 459.820000 83.840000 ;
      RECT 371.620000 82.760000 414.820000 83.840000 ;
      RECT 326.620000 82.760000 369.820000 83.840000 ;
      RECT 281.620000 82.760000 324.820000 83.840000 ;
      RECT 236.620000 82.760000 279.820000 83.840000 ;
      RECT 191.620000 82.760000 234.820000 83.840000 ;
      RECT 146.620000 82.760000 189.820000 83.840000 ;
      RECT 101.620000 82.760000 144.820000 83.840000 ;
      RECT 56.620000 82.760000 99.820000 83.840000 ;
      RECT 11.620000 82.760000 54.820000 83.840000 ;
      RECT 4.860000 82.760000 9.655000 83.840000 ;
      RECT 0.000000 82.760000 3.060000 83.840000 ;
      RECT 0.000000 82.500000 550.160000 82.760000 ;
      RECT 0.000000 81.520000 548.960000 82.500000 ;
      RECT 0.000000 81.120000 550.160000 81.520000 ;
      RECT 544.900000 80.040000 550.160000 81.120000 ;
      RECT 508.620000 80.040000 543.100000 81.120000 ;
      RECT 463.620000 80.040000 506.820000 81.120000 ;
      RECT 418.620000 80.040000 461.820000 81.120000 ;
      RECT 373.620000 80.040000 416.820000 81.120000 ;
      RECT 328.620000 80.040000 371.820000 81.120000 ;
      RECT 283.620000 80.040000 326.820000 81.120000 ;
      RECT 238.620000 80.040000 281.820000 81.120000 ;
      RECT 193.620000 80.040000 236.820000 81.120000 ;
      RECT 148.620000 80.040000 191.820000 81.120000 ;
      RECT 103.620000 80.040000 146.820000 81.120000 ;
      RECT 58.620000 80.040000 101.820000 81.120000 ;
      RECT 13.620000 80.040000 56.820000 81.120000 ;
      RECT 7.060000 80.040000 11.820000 81.120000 ;
      RECT 0.000000 80.040000 5.260000 81.120000 ;
      RECT 0.000000 79.450000 550.160000 80.040000 ;
      RECT 0.000000 78.470000 548.960000 79.450000 ;
      RECT 0.000000 78.400000 550.160000 78.470000 ;
      RECT 547.100000 77.320000 550.160000 78.400000 ;
      RECT 506.620000 77.320000 545.300000 78.400000 ;
      RECT 461.620000 77.320000 504.820000 78.400000 ;
      RECT 416.620000 77.320000 459.820000 78.400000 ;
      RECT 371.620000 77.320000 414.820000 78.400000 ;
      RECT 326.620000 77.320000 369.820000 78.400000 ;
      RECT 281.620000 77.320000 324.820000 78.400000 ;
      RECT 236.620000 77.320000 279.820000 78.400000 ;
      RECT 191.620000 77.320000 234.820000 78.400000 ;
      RECT 146.620000 77.320000 189.820000 78.400000 ;
      RECT 101.620000 77.320000 144.820000 78.400000 ;
      RECT 56.620000 77.320000 99.820000 78.400000 ;
      RECT 11.620000 77.320000 54.820000 78.400000 ;
      RECT 4.860000 77.320000 9.655000 78.400000 ;
      RECT 0.000000 77.320000 3.060000 78.400000 ;
      RECT 0.000000 75.790000 550.160000 77.320000 ;
      RECT 0.000000 75.680000 548.960000 75.790000 ;
      RECT 544.900000 74.810000 548.960000 75.680000 ;
      RECT 544.900000 74.600000 550.160000 74.810000 ;
      RECT 508.620000 74.600000 543.100000 75.680000 ;
      RECT 463.620000 74.600000 506.820000 75.680000 ;
      RECT 418.620000 74.600000 461.820000 75.680000 ;
      RECT 373.620000 74.600000 416.820000 75.680000 ;
      RECT 328.620000 74.600000 371.820000 75.680000 ;
      RECT 283.620000 74.600000 326.820000 75.680000 ;
      RECT 238.620000 74.600000 281.820000 75.680000 ;
      RECT 193.620000 74.600000 236.820000 75.680000 ;
      RECT 148.620000 74.600000 191.820000 75.680000 ;
      RECT 103.620000 74.600000 146.820000 75.680000 ;
      RECT 58.620000 74.600000 101.820000 75.680000 ;
      RECT 13.620000 74.600000 56.820000 75.680000 ;
      RECT 7.060000 74.600000 11.820000 75.680000 ;
      RECT 0.000000 74.600000 5.260000 75.680000 ;
      RECT 0.000000 72.960000 550.160000 74.600000 ;
      RECT 547.100000 72.130000 550.160000 72.960000 ;
      RECT 547.100000 71.880000 548.960000 72.130000 ;
      RECT 506.620000 71.880000 545.300000 72.960000 ;
      RECT 461.620000 71.880000 504.820000 72.960000 ;
      RECT 416.620000 71.880000 459.820000 72.960000 ;
      RECT 371.620000 71.880000 414.820000 72.960000 ;
      RECT 326.620000 71.880000 369.820000 72.960000 ;
      RECT 281.620000 71.880000 324.820000 72.960000 ;
      RECT 236.620000 71.880000 279.820000 72.960000 ;
      RECT 191.620000 71.880000 234.820000 72.960000 ;
      RECT 146.620000 71.880000 189.820000 72.960000 ;
      RECT 101.620000 71.880000 144.820000 72.960000 ;
      RECT 56.620000 71.880000 99.820000 72.960000 ;
      RECT 11.620000 71.880000 54.820000 72.960000 ;
      RECT 4.860000 71.880000 9.655000 72.960000 ;
      RECT 0.000000 71.880000 3.060000 72.960000 ;
      RECT 0.000000 71.150000 548.960000 71.880000 ;
      RECT 0.000000 70.240000 550.160000 71.150000 ;
      RECT 544.900000 69.160000 550.160000 70.240000 ;
      RECT 508.620000 69.160000 543.100000 70.240000 ;
      RECT 463.620000 69.160000 506.820000 70.240000 ;
      RECT 418.620000 69.160000 461.820000 70.240000 ;
      RECT 373.620000 69.160000 416.820000 70.240000 ;
      RECT 328.620000 69.160000 371.820000 70.240000 ;
      RECT 283.620000 69.160000 326.820000 70.240000 ;
      RECT 238.620000 69.160000 281.820000 70.240000 ;
      RECT 193.620000 69.160000 236.820000 70.240000 ;
      RECT 148.620000 69.160000 191.820000 70.240000 ;
      RECT 103.620000 69.160000 146.820000 70.240000 ;
      RECT 58.620000 69.160000 101.820000 70.240000 ;
      RECT 13.620000 69.160000 56.820000 70.240000 ;
      RECT 7.060000 69.160000 11.820000 70.240000 ;
      RECT 0.000000 69.160000 5.260000 70.240000 ;
      RECT 0.000000 69.080000 550.160000 69.160000 ;
      RECT 0.000000 68.100000 548.960000 69.080000 ;
      RECT 0.000000 67.520000 550.160000 68.100000 ;
      RECT 547.100000 66.440000 550.160000 67.520000 ;
      RECT 506.620000 66.440000 545.300000 67.520000 ;
      RECT 461.620000 66.440000 504.820000 67.520000 ;
      RECT 416.620000 66.440000 459.820000 67.520000 ;
      RECT 371.620000 66.440000 414.820000 67.520000 ;
      RECT 326.620000 66.440000 369.820000 67.520000 ;
      RECT 281.620000 66.440000 324.820000 67.520000 ;
      RECT 236.620000 66.440000 279.820000 67.520000 ;
      RECT 191.620000 66.440000 234.820000 67.520000 ;
      RECT 146.620000 66.440000 189.820000 67.520000 ;
      RECT 101.620000 66.440000 144.820000 67.520000 ;
      RECT 56.620000 66.440000 99.820000 67.520000 ;
      RECT 11.620000 66.440000 54.820000 67.520000 ;
      RECT 4.860000 66.440000 9.655000 67.520000 ;
      RECT 0.000000 66.440000 3.060000 67.520000 ;
      RECT 0.000000 65.420000 550.160000 66.440000 ;
      RECT 0.000000 64.800000 548.960000 65.420000 ;
      RECT 544.900000 64.440000 548.960000 64.800000 ;
      RECT 544.900000 63.720000 550.160000 64.440000 ;
      RECT 508.620000 63.720000 543.100000 64.800000 ;
      RECT 463.620000 63.720000 506.820000 64.800000 ;
      RECT 418.620000 63.720000 461.820000 64.800000 ;
      RECT 373.620000 63.720000 416.820000 64.800000 ;
      RECT 328.620000 63.720000 371.820000 64.800000 ;
      RECT 283.620000 63.720000 326.820000 64.800000 ;
      RECT 238.620000 63.720000 281.820000 64.800000 ;
      RECT 193.620000 63.720000 236.820000 64.800000 ;
      RECT 148.620000 63.720000 191.820000 64.800000 ;
      RECT 103.620000 63.720000 146.820000 64.800000 ;
      RECT 58.620000 63.720000 101.820000 64.800000 ;
      RECT 13.620000 63.720000 56.820000 64.800000 ;
      RECT 7.060000 63.720000 11.820000 64.800000 ;
      RECT 0.000000 63.720000 5.260000 64.800000 ;
      RECT 0.000000 62.080000 550.160000 63.720000 ;
      RECT 547.100000 61.760000 550.160000 62.080000 ;
      RECT 547.100000 61.000000 548.960000 61.760000 ;
      RECT 506.620000 61.000000 545.300000 62.080000 ;
      RECT 461.620000 61.000000 504.820000 62.080000 ;
      RECT 416.620000 61.000000 459.820000 62.080000 ;
      RECT 371.620000 61.000000 414.820000 62.080000 ;
      RECT 326.620000 61.000000 369.820000 62.080000 ;
      RECT 281.620000 61.000000 324.820000 62.080000 ;
      RECT 236.620000 61.000000 279.820000 62.080000 ;
      RECT 191.620000 61.000000 234.820000 62.080000 ;
      RECT 146.620000 61.000000 189.820000 62.080000 ;
      RECT 101.620000 61.000000 144.820000 62.080000 ;
      RECT 56.620000 61.000000 99.820000 62.080000 ;
      RECT 11.620000 61.000000 54.820000 62.080000 ;
      RECT 4.860000 61.000000 9.655000 62.080000 ;
      RECT 0.000000 61.000000 3.060000 62.080000 ;
      RECT 0.000000 60.780000 548.960000 61.000000 ;
      RECT 0.000000 59.360000 550.160000 60.780000 ;
      RECT 544.900000 58.710000 550.160000 59.360000 ;
      RECT 544.900000 58.280000 548.960000 58.710000 ;
      RECT 508.620000 58.280000 543.100000 59.360000 ;
      RECT 463.620000 58.280000 506.820000 59.360000 ;
      RECT 418.620000 58.280000 461.820000 59.360000 ;
      RECT 373.620000 58.280000 416.820000 59.360000 ;
      RECT 328.620000 58.280000 371.820000 59.360000 ;
      RECT 283.620000 58.280000 326.820000 59.360000 ;
      RECT 238.620000 58.280000 281.820000 59.360000 ;
      RECT 193.620000 58.280000 236.820000 59.360000 ;
      RECT 148.620000 58.280000 191.820000 59.360000 ;
      RECT 103.620000 58.280000 146.820000 59.360000 ;
      RECT 58.620000 58.280000 101.820000 59.360000 ;
      RECT 13.620000 58.280000 56.820000 59.360000 ;
      RECT 7.060000 58.280000 11.820000 59.360000 ;
      RECT 0.000000 58.280000 5.260000 59.360000 ;
      RECT 0.000000 57.730000 548.960000 58.280000 ;
      RECT 0.000000 56.640000 550.160000 57.730000 ;
      RECT 547.100000 55.560000 550.160000 56.640000 ;
      RECT 506.620000 55.560000 545.300000 56.640000 ;
      RECT 461.620000 55.560000 504.820000 56.640000 ;
      RECT 416.620000 55.560000 459.820000 56.640000 ;
      RECT 371.620000 55.560000 414.820000 56.640000 ;
      RECT 326.620000 55.560000 369.820000 56.640000 ;
      RECT 281.620000 55.560000 324.820000 56.640000 ;
      RECT 236.620000 55.560000 279.820000 56.640000 ;
      RECT 191.620000 55.560000 234.820000 56.640000 ;
      RECT 146.620000 55.560000 189.820000 56.640000 ;
      RECT 101.620000 55.560000 144.820000 56.640000 ;
      RECT 56.620000 55.560000 99.820000 56.640000 ;
      RECT 11.620000 55.560000 54.820000 56.640000 ;
      RECT 4.860000 55.560000 9.655000 56.640000 ;
      RECT 0.000000 55.560000 3.060000 56.640000 ;
      RECT 0.000000 55.050000 550.160000 55.560000 ;
      RECT 0.000000 54.070000 548.960000 55.050000 ;
      RECT 0.000000 53.920000 550.160000 54.070000 ;
      RECT 544.900000 52.840000 550.160000 53.920000 ;
      RECT 508.620000 52.840000 543.100000 53.920000 ;
      RECT 463.620000 52.840000 506.820000 53.920000 ;
      RECT 418.620000 52.840000 461.820000 53.920000 ;
      RECT 373.620000 52.840000 416.820000 53.920000 ;
      RECT 328.620000 52.840000 371.820000 53.920000 ;
      RECT 283.620000 52.840000 326.820000 53.920000 ;
      RECT 238.620000 52.840000 281.820000 53.920000 ;
      RECT 193.620000 52.840000 236.820000 53.920000 ;
      RECT 148.620000 52.840000 191.820000 53.920000 ;
      RECT 103.620000 52.840000 146.820000 53.920000 ;
      RECT 58.620000 52.840000 101.820000 53.920000 ;
      RECT 13.620000 52.840000 56.820000 53.920000 ;
      RECT 7.060000 52.840000 11.820000 53.920000 ;
      RECT 0.000000 52.840000 5.260000 53.920000 ;
      RECT 0.000000 51.390000 550.160000 52.840000 ;
      RECT 0.000000 51.200000 548.960000 51.390000 ;
      RECT 547.100000 50.410000 548.960000 51.200000 ;
      RECT 547.100000 50.120000 550.160000 50.410000 ;
      RECT 506.620000 50.120000 545.300000 51.200000 ;
      RECT 461.620000 50.120000 504.820000 51.200000 ;
      RECT 416.620000 50.120000 459.820000 51.200000 ;
      RECT 371.620000 50.120000 414.820000 51.200000 ;
      RECT 326.620000 50.120000 369.820000 51.200000 ;
      RECT 281.620000 50.120000 324.820000 51.200000 ;
      RECT 236.620000 50.120000 279.820000 51.200000 ;
      RECT 191.620000 50.120000 234.820000 51.200000 ;
      RECT 146.620000 50.120000 189.820000 51.200000 ;
      RECT 101.620000 50.120000 144.820000 51.200000 ;
      RECT 56.620000 50.120000 99.820000 51.200000 ;
      RECT 11.620000 50.120000 54.820000 51.200000 ;
      RECT 4.860000 50.120000 9.655000 51.200000 ;
      RECT 0.000000 50.120000 3.060000 51.200000 ;
      RECT 0.000000 48.480000 550.160000 50.120000 ;
      RECT 544.900000 48.340000 550.160000 48.480000 ;
      RECT 544.900000 47.400000 548.960000 48.340000 ;
      RECT 508.620000 47.400000 543.100000 48.480000 ;
      RECT 463.620000 47.400000 506.820000 48.480000 ;
      RECT 418.620000 47.400000 461.820000 48.480000 ;
      RECT 373.620000 47.400000 416.820000 48.480000 ;
      RECT 328.620000 47.400000 371.820000 48.480000 ;
      RECT 283.620000 47.400000 326.820000 48.480000 ;
      RECT 238.620000 47.400000 281.820000 48.480000 ;
      RECT 193.620000 47.400000 236.820000 48.480000 ;
      RECT 148.620000 47.400000 191.820000 48.480000 ;
      RECT 103.620000 47.400000 146.820000 48.480000 ;
      RECT 58.620000 47.400000 101.820000 48.480000 ;
      RECT 13.620000 47.400000 56.820000 48.480000 ;
      RECT 7.060000 47.400000 11.820000 48.480000 ;
      RECT 0.000000 47.400000 5.260000 48.480000 ;
      RECT 0.000000 47.360000 548.960000 47.400000 ;
      RECT 0.000000 45.760000 550.160000 47.360000 ;
      RECT 547.100000 44.680000 550.160000 45.760000 ;
      RECT 506.620000 44.680000 545.300000 45.760000 ;
      RECT 461.620000 44.680000 504.820000 45.760000 ;
      RECT 416.620000 44.680000 459.820000 45.760000 ;
      RECT 371.620000 44.680000 414.820000 45.760000 ;
      RECT 326.620000 44.680000 369.820000 45.760000 ;
      RECT 281.620000 44.680000 324.820000 45.760000 ;
      RECT 236.620000 44.680000 279.820000 45.760000 ;
      RECT 191.620000 44.680000 234.820000 45.760000 ;
      RECT 146.620000 44.680000 189.820000 45.760000 ;
      RECT 101.620000 44.680000 144.820000 45.760000 ;
      RECT 56.620000 44.680000 99.820000 45.760000 ;
      RECT 11.620000 44.680000 54.820000 45.760000 ;
      RECT 4.860000 44.680000 9.655000 45.760000 ;
      RECT 0.000000 44.680000 3.060000 45.760000 ;
      RECT 0.000000 43.700000 548.960000 44.680000 ;
      RECT 0.000000 43.040000 550.160000 43.700000 ;
      RECT 544.900000 41.960000 550.160000 43.040000 ;
      RECT 508.620000 41.960000 543.100000 43.040000 ;
      RECT 463.620000 41.960000 506.820000 43.040000 ;
      RECT 418.620000 41.960000 461.820000 43.040000 ;
      RECT 373.620000 41.960000 416.820000 43.040000 ;
      RECT 328.620000 41.960000 371.820000 43.040000 ;
      RECT 283.620000 41.960000 326.820000 43.040000 ;
      RECT 238.620000 41.960000 281.820000 43.040000 ;
      RECT 193.620000 41.960000 236.820000 43.040000 ;
      RECT 148.620000 41.960000 191.820000 43.040000 ;
      RECT 103.620000 41.960000 146.820000 43.040000 ;
      RECT 58.620000 41.960000 101.820000 43.040000 ;
      RECT 13.620000 41.960000 56.820000 43.040000 ;
      RECT 7.060000 41.960000 11.820000 43.040000 ;
      RECT 0.000000 41.960000 5.260000 43.040000 ;
      RECT 0.000000 41.020000 550.160000 41.960000 ;
      RECT 0.000000 40.320000 548.960000 41.020000 ;
      RECT 547.100000 40.040000 548.960000 40.320000 ;
      RECT 547.100000 39.240000 550.160000 40.040000 ;
      RECT 506.620000 39.240000 545.300000 40.320000 ;
      RECT 461.620000 39.240000 504.820000 40.320000 ;
      RECT 416.620000 39.240000 459.820000 40.320000 ;
      RECT 371.620000 39.240000 414.820000 40.320000 ;
      RECT 326.620000 39.240000 369.820000 40.320000 ;
      RECT 281.620000 39.240000 324.820000 40.320000 ;
      RECT 236.620000 39.240000 279.820000 40.320000 ;
      RECT 191.620000 39.240000 234.820000 40.320000 ;
      RECT 146.620000 39.240000 189.820000 40.320000 ;
      RECT 101.620000 39.240000 144.820000 40.320000 ;
      RECT 56.620000 39.240000 99.820000 40.320000 ;
      RECT 11.620000 39.240000 54.820000 40.320000 ;
      RECT 4.860000 39.240000 9.655000 40.320000 ;
      RECT 0.000000 39.240000 3.060000 40.320000 ;
      RECT 0.000000 37.970000 550.160000 39.240000 ;
      RECT 0.000000 37.600000 548.960000 37.970000 ;
      RECT 544.900000 36.990000 548.960000 37.600000 ;
      RECT 544.900000 36.520000 550.160000 36.990000 ;
      RECT 508.620000 36.520000 543.100000 37.600000 ;
      RECT 463.620000 36.520000 506.820000 37.600000 ;
      RECT 418.620000 36.520000 461.820000 37.600000 ;
      RECT 373.620000 36.520000 416.820000 37.600000 ;
      RECT 328.620000 36.520000 371.820000 37.600000 ;
      RECT 283.620000 36.520000 326.820000 37.600000 ;
      RECT 238.620000 36.520000 281.820000 37.600000 ;
      RECT 193.620000 36.520000 236.820000 37.600000 ;
      RECT 148.620000 36.520000 191.820000 37.600000 ;
      RECT 103.620000 36.520000 146.820000 37.600000 ;
      RECT 58.620000 36.520000 101.820000 37.600000 ;
      RECT 13.620000 36.520000 56.820000 37.600000 ;
      RECT 7.060000 36.520000 11.820000 37.600000 ;
      RECT 0.000000 36.520000 5.260000 37.600000 ;
      RECT 0.000000 34.880000 550.160000 36.520000 ;
      RECT 547.100000 34.310000 550.160000 34.880000 ;
      RECT 547.100000 33.800000 548.960000 34.310000 ;
      RECT 506.620000 33.800000 545.300000 34.880000 ;
      RECT 461.620000 33.800000 504.820000 34.880000 ;
      RECT 416.620000 33.800000 459.820000 34.880000 ;
      RECT 371.620000 33.800000 414.820000 34.880000 ;
      RECT 326.620000 33.800000 369.820000 34.880000 ;
      RECT 281.620000 33.800000 324.820000 34.880000 ;
      RECT 236.620000 33.800000 279.820000 34.880000 ;
      RECT 191.620000 33.800000 234.820000 34.880000 ;
      RECT 146.620000 33.800000 189.820000 34.880000 ;
      RECT 101.620000 33.800000 144.820000 34.880000 ;
      RECT 56.620000 33.800000 99.820000 34.880000 ;
      RECT 11.620000 33.800000 54.820000 34.880000 ;
      RECT 4.860000 33.800000 9.655000 34.880000 ;
      RECT 0.000000 33.800000 3.060000 34.880000 ;
      RECT 0.000000 33.330000 548.960000 33.800000 ;
      RECT 0.000000 32.160000 550.160000 33.330000 ;
      RECT 544.900000 31.080000 550.160000 32.160000 ;
      RECT 508.620000 31.080000 543.100000 32.160000 ;
      RECT 463.620000 31.080000 506.820000 32.160000 ;
      RECT 418.620000 31.080000 461.820000 32.160000 ;
      RECT 373.620000 31.080000 416.820000 32.160000 ;
      RECT 328.620000 31.080000 371.820000 32.160000 ;
      RECT 283.620000 31.080000 326.820000 32.160000 ;
      RECT 238.620000 31.080000 281.820000 32.160000 ;
      RECT 193.620000 31.080000 236.820000 32.160000 ;
      RECT 148.620000 31.080000 191.820000 32.160000 ;
      RECT 103.620000 31.080000 146.820000 32.160000 ;
      RECT 58.620000 31.080000 101.820000 32.160000 ;
      RECT 13.620000 31.080000 56.820000 32.160000 ;
      RECT 7.060000 31.080000 11.820000 32.160000 ;
      RECT 0.000000 31.080000 5.260000 32.160000 ;
      RECT 0.000000 30.650000 550.160000 31.080000 ;
      RECT 0.000000 29.670000 548.960000 30.650000 ;
      RECT 0.000000 29.440000 550.160000 29.670000 ;
      RECT 547.100000 28.360000 550.160000 29.440000 ;
      RECT 506.620000 28.360000 545.300000 29.440000 ;
      RECT 461.620000 28.360000 504.820000 29.440000 ;
      RECT 416.620000 28.360000 459.820000 29.440000 ;
      RECT 371.620000 28.360000 414.820000 29.440000 ;
      RECT 326.620000 28.360000 369.820000 29.440000 ;
      RECT 281.620000 28.360000 324.820000 29.440000 ;
      RECT 236.620000 28.360000 279.820000 29.440000 ;
      RECT 191.620000 28.360000 234.820000 29.440000 ;
      RECT 146.620000 28.360000 189.820000 29.440000 ;
      RECT 101.620000 28.360000 144.820000 29.440000 ;
      RECT 56.620000 28.360000 99.820000 29.440000 ;
      RECT 11.620000 28.360000 54.820000 29.440000 ;
      RECT 4.860000 28.360000 9.655000 29.440000 ;
      RECT 0.000000 28.360000 3.060000 29.440000 ;
      RECT 0.000000 27.600000 550.160000 28.360000 ;
      RECT 0.000000 26.720000 548.960000 27.600000 ;
      RECT 544.900000 26.620000 548.960000 26.720000 ;
      RECT 544.900000 25.640000 550.160000 26.620000 ;
      RECT 508.620000 25.640000 543.100000 26.720000 ;
      RECT 463.620000 25.640000 506.820000 26.720000 ;
      RECT 418.620000 25.640000 461.820000 26.720000 ;
      RECT 373.620000 25.640000 416.820000 26.720000 ;
      RECT 328.620000 25.640000 371.820000 26.720000 ;
      RECT 283.620000 25.640000 326.820000 26.720000 ;
      RECT 238.620000 25.640000 281.820000 26.720000 ;
      RECT 193.620000 25.640000 236.820000 26.720000 ;
      RECT 148.620000 25.640000 191.820000 26.720000 ;
      RECT 103.620000 25.640000 146.820000 26.720000 ;
      RECT 58.620000 25.640000 101.820000 26.720000 ;
      RECT 13.620000 25.640000 56.820000 26.720000 ;
      RECT 7.060000 25.640000 11.820000 26.720000 ;
      RECT 0.000000 25.640000 5.260000 26.720000 ;
      RECT 0.000000 24.000000 550.160000 25.640000 ;
      RECT 547.100000 23.940000 550.160000 24.000000 ;
      RECT 547.100000 22.960000 548.960000 23.940000 ;
      RECT 547.100000 22.920000 550.160000 22.960000 ;
      RECT 506.620000 22.920000 545.300000 24.000000 ;
      RECT 461.620000 22.920000 504.820000 24.000000 ;
      RECT 416.620000 22.920000 459.820000 24.000000 ;
      RECT 371.620000 22.920000 414.820000 24.000000 ;
      RECT 326.620000 22.920000 369.820000 24.000000 ;
      RECT 281.620000 22.920000 324.820000 24.000000 ;
      RECT 236.620000 22.920000 279.820000 24.000000 ;
      RECT 191.620000 22.920000 234.820000 24.000000 ;
      RECT 146.620000 22.920000 189.820000 24.000000 ;
      RECT 101.620000 22.920000 144.820000 24.000000 ;
      RECT 56.620000 22.920000 99.820000 24.000000 ;
      RECT 11.620000 22.920000 54.820000 24.000000 ;
      RECT 4.860000 22.920000 9.655000 24.000000 ;
      RECT 0.000000 22.920000 3.060000 24.000000 ;
      RECT 0.000000 21.280000 550.160000 22.920000 ;
      RECT 544.900000 20.280000 550.160000 21.280000 ;
      RECT 544.900000 20.200000 548.960000 20.280000 ;
      RECT 508.620000 20.200000 543.100000 21.280000 ;
      RECT 463.620000 20.200000 506.820000 21.280000 ;
      RECT 418.620000 20.200000 461.820000 21.280000 ;
      RECT 373.620000 20.200000 416.820000 21.280000 ;
      RECT 328.620000 20.200000 371.820000 21.280000 ;
      RECT 283.620000 20.200000 326.820000 21.280000 ;
      RECT 238.620000 20.200000 281.820000 21.280000 ;
      RECT 193.620000 20.200000 236.820000 21.280000 ;
      RECT 148.620000 20.200000 191.820000 21.280000 ;
      RECT 103.620000 20.200000 146.820000 21.280000 ;
      RECT 58.620000 20.200000 101.820000 21.280000 ;
      RECT 13.620000 20.200000 56.820000 21.280000 ;
      RECT 7.060000 20.200000 11.820000 21.280000 ;
      RECT 0.000000 20.200000 5.260000 21.280000 ;
      RECT 0.000000 19.300000 548.960000 20.200000 ;
      RECT 0.000000 18.560000 550.160000 19.300000 ;
      RECT 547.100000 17.480000 550.160000 18.560000 ;
      RECT 506.620000 17.480000 545.300000 18.560000 ;
      RECT 461.620000 17.480000 504.820000 18.560000 ;
      RECT 416.620000 17.480000 459.820000 18.560000 ;
      RECT 371.620000 17.480000 414.820000 18.560000 ;
      RECT 326.620000 17.480000 369.820000 18.560000 ;
      RECT 281.620000 17.480000 324.820000 18.560000 ;
      RECT 236.620000 17.480000 279.820000 18.560000 ;
      RECT 191.620000 17.480000 234.820000 18.560000 ;
      RECT 146.620000 17.480000 189.820000 18.560000 ;
      RECT 101.620000 17.480000 144.820000 18.560000 ;
      RECT 56.620000 17.480000 99.820000 18.560000 ;
      RECT 11.620000 17.480000 54.820000 18.560000 ;
      RECT 4.860000 17.480000 9.655000 18.560000 ;
      RECT 0.000000 17.480000 3.060000 18.560000 ;
      RECT 0.000000 17.230000 550.160000 17.480000 ;
      RECT 0.000000 16.250000 548.960000 17.230000 ;
      RECT 0.000000 15.840000 550.160000 16.250000 ;
      RECT 544.900000 14.760000 550.160000 15.840000 ;
      RECT 508.620000 14.760000 543.100000 15.840000 ;
      RECT 463.620000 14.760000 506.820000 15.840000 ;
      RECT 418.620000 14.760000 461.820000 15.840000 ;
      RECT 373.620000 14.760000 416.820000 15.840000 ;
      RECT 328.620000 14.760000 371.820000 15.840000 ;
      RECT 283.620000 14.760000 326.820000 15.840000 ;
      RECT 238.620000 14.760000 281.820000 15.840000 ;
      RECT 193.620000 14.760000 236.820000 15.840000 ;
      RECT 148.620000 14.760000 191.820000 15.840000 ;
      RECT 103.620000 14.760000 146.820000 15.840000 ;
      RECT 58.620000 14.760000 101.820000 15.840000 ;
      RECT 13.620000 14.760000 56.820000 15.840000 ;
      RECT 7.060000 14.760000 11.820000 15.840000 ;
      RECT 0.000000 14.760000 5.260000 15.840000 ;
      RECT 0.000000 13.570000 550.160000 14.760000 ;
      RECT 0.000000 13.120000 548.960000 13.570000 ;
      RECT 547.100000 12.590000 548.960000 13.120000 ;
      RECT 547.100000 12.040000 550.160000 12.590000 ;
      RECT 506.620000 12.040000 545.300000 13.120000 ;
      RECT 461.620000 12.040000 504.820000 13.120000 ;
      RECT 416.620000 12.040000 459.820000 13.120000 ;
      RECT 371.620000 12.040000 414.820000 13.120000 ;
      RECT 326.620000 12.040000 369.820000 13.120000 ;
      RECT 281.620000 12.040000 324.820000 13.120000 ;
      RECT 236.620000 12.040000 279.820000 13.120000 ;
      RECT 191.620000 12.040000 234.820000 13.120000 ;
      RECT 146.620000 12.040000 189.820000 13.120000 ;
      RECT 101.620000 12.040000 144.820000 13.120000 ;
      RECT 56.620000 12.040000 99.820000 13.120000 ;
      RECT 11.620000 12.040000 54.820000 13.120000 ;
      RECT 4.860000 12.040000 9.655000 13.120000 ;
      RECT 0.000000 12.040000 3.060000 13.120000 ;
      RECT 0.000000 10.520000 550.160000 12.040000 ;
      RECT 0.000000 10.400000 548.960000 10.520000 ;
      RECT 544.900000 9.540000 548.960000 10.400000 ;
      RECT 544.900000 9.320000 550.160000 9.540000 ;
      RECT 508.620000 9.320000 543.100000 10.400000 ;
      RECT 463.620000 9.320000 506.820000 10.400000 ;
      RECT 418.620000 9.320000 461.820000 10.400000 ;
      RECT 373.620000 9.320000 416.820000 10.400000 ;
      RECT 328.620000 9.320000 371.820000 10.400000 ;
      RECT 283.620000 9.320000 326.820000 10.400000 ;
      RECT 238.620000 9.320000 281.820000 10.400000 ;
      RECT 193.620000 9.320000 236.820000 10.400000 ;
      RECT 148.620000 9.320000 191.820000 10.400000 ;
      RECT 103.620000 9.320000 146.820000 10.400000 ;
      RECT 58.620000 9.320000 101.820000 10.400000 ;
      RECT 13.620000 9.320000 56.820000 10.400000 ;
      RECT 7.060000 9.320000 11.820000 10.400000 ;
      RECT 0.000000 9.320000 5.260000 10.400000 ;
      RECT 0.000000 6.930000 550.160000 9.320000 ;
      RECT 0.000000 4.730000 550.160000 5.130000 ;
      RECT 0.000000 0.000000 550.160000 2.930000 ;
    LAYER met4 ;
      RECT 7.060000 596.490000 543.100000 599.760000 ;
      RECT 506.620000 594.290000 543.100000 596.490000 ;
      RECT 461.620000 594.290000 504.820000 596.490000 ;
      RECT 416.620000 594.290000 459.820000 596.490000 ;
      RECT 371.620000 594.290000 414.820000 596.490000 ;
      RECT 326.620000 594.290000 369.820000 596.490000 ;
      RECT 281.620000 594.290000 324.820000 596.490000 ;
      RECT 236.620000 594.290000 279.820000 596.490000 ;
      RECT 191.620000 594.290000 234.820000 596.490000 ;
      RECT 146.620000 594.290000 189.820000 596.490000 ;
      RECT 101.620000 594.290000 144.820000 596.490000 ;
      RECT 56.620000 594.290000 99.820000 596.490000 ;
      RECT 11.620000 594.290000 54.820000 596.490000 ;
      RECT 7.060000 589.760000 9.820000 596.490000 ;
      RECT 7.060000 588.680000 9.655000 589.760000 ;
      RECT 7.060000 584.320000 9.820000 588.680000 ;
      RECT 7.060000 583.240000 9.655000 584.320000 ;
      RECT 7.060000 578.880000 9.820000 583.240000 ;
      RECT 7.060000 577.800000 9.655000 578.880000 ;
      RECT 7.060000 573.440000 9.820000 577.800000 ;
      RECT 7.060000 572.360000 9.655000 573.440000 ;
      RECT 7.060000 568.000000 9.820000 572.360000 ;
      RECT 7.060000 566.920000 9.655000 568.000000 ;
      RECT 7.060000 562.560000 9.820000 566.920000 ;
      RECT 7.060000 561.480000 9.655000 562.560000 ;
      RECT 7.060000 557.120000 9.820000 561.480000 ;
      RECT 7.060000 556.040000 9.655000 557.120000 ;
      RECT 7.060000 551.680000 9.820000 556.040000 ;
      RECT 7.060000 550.600000 9.655000 551.680000 ;
      RECT 7.060000 546.240000 9.820000 550.600000 ;
      RECT 7.060000 545.160000 9.655000 546.240000 ;
      RECT 7.060000 540.800000 9.820000 545.160000 ;
      RECT 7.060000 539.720000 9.655000 540.800000 ;
      RECT 7.060000 535.360000 9.820000 539.720000 ;
      RECT 7.060000 534.280000 9.655000 535.360000 ;
      RECT 7.060000 529.920000 9.820000 534.280000 ;
      RECT 7.060000 528.840000 9.655000 529.920000 ;
      RECT 7.060000 524.480000 9.820000 528.840000 ;
      RECT 7.060000 523.400000 9.655000 524.480000 ;
      RECT 7.060000 519.040000 9.820000 523.400000 ;
      RECT 7.060000 517.960000 9.655000 519.040000 ;
      RECT 7.060000 513.600000 9.820000 517.960000 ;
      RECT 7.060000 512.520000 9.655000 513.600000 ;
      RECT 7.060000 508.160000 9.820000 512.520000 ;
      RECT 7.060000 507.080000 9.655000 508.160000 ;
      RECT 7.060000 502.720000 9.820000 507.080000 ;
      RECT 7.060000 501.640000 9.655000 502.720000 ;
      RECT 7.060000 497.280000 9.820000 501.640000 ;
      RECT 7.060000 496.200000 9.655000 497.280000 ;
      RECT 7.060000 491.840000 9.820000 496.200000 ;
      RECT 7.060000 490.760000 9.655000 491.840000 ;
      RECT 7.060000 486.400000 9.820000 490.760000 ;
      RECT 7.060000 485.320000 9.655000 486.400000 ;
      RECT 7.060000 480.960000 9.820000 485.320000 ;
      RECT 7.060000 479.880000 9.655000 480.960000 ;
      RECT 7.060000 475.520000 9.820000 479.880000 ;
      RECT 7.060000 474.440000 9.655000 475.520000 ;
      RECT 7.060000 470.080000 9.820000 474.440000 ;
      RECT 7.060000 469.000000 9.655000 470.080000 ;
      RECT 7.060000 464.640000 9.820000 469.000000 ;
      RECT 7.060000 463.560000 9.655000 464.640000 ;
      RECT 7.060000 459.200000 9.820000 463.560000 ;
      RECT 7.060000 458.120000 9.655000 459.200000 ;
      RECT 7.060000 453.760000 9.820000 458.120000 ;
      RECT 7.060000 452.680000 9.655000 453.760000 ;
      RECT 7.060000 448.320000 9.820000 452.680000 ;
      RECT 7.060000 447.240000 9.655000 448.320000 ;
      RECT 7.060000 442.880000 9.820000 447.240000 ;
      RECT 7.060000 441.800000 9.655000 442.880000 ;
      RECT 7.060000 437.440000 9.820000 441.800000 ;
      RECT 7.060000 436.360000 9.655000 437.440000 ;
      RECT 7.060000 432.000000 9.820000 436.360000 ;
      RECT 7.060000 430.920000 9.655000 432.000000 ;
      RECT 7.060000 426.560000 9.820000 430.920000 ;
      RECT 7.060000 425.480000 9.655000 426.560000 ;
      RECT 7.060000 421.120000 9.820000 425.480000 ;
      RECT 7.060000 420.040000 9.655000 421.120000 ;
      RECT 7.060000 415.680000 9.820000 420.040000 ;
      RECT 7.060000 414.600000 9.655000 415.680000 ;
      RECT 7.060000 410.240000 9.820000 414.600000 ;
      RECT 7.060000 409.160000 9.655000 410.240000 ;
      RECT 7.060000 404.800000 9.820000 409.160000 ;
      RECT 7.060000 403.720000 9.655000 404.800000 ;
      RECT 7.060000 399.360000 9.820000 403.720000 ;
      RECT 7.060000 398.280000 9.655000 399.360000 ;
      RECT 7.060000 393.920000 9.820000 398.280000 ;
      RECT 7.060000 392.840000 9.655000 393.920000 ;
      RECT 7.060000 388.480000 9.820000 392.840000 ;
      RECT 7.060000 387.400000 9.655000 388.480000 ;
      RECT 7.060000 383.040000 9.820000 387.400000 ;
      RECT 7.060000 381.960000 9.655000 383.040000 ;
      RECT 7.060000 377.600000 9.820000 381.960000 ;
      RECT 7.060000 376.520000 9.655000 377.600000 ;
      RECT 7.060000 372.160000 9.820000 376.520000 ;
      RECT 7.060000 371.080000 9.655000 372.160000 ;
      RECT 7.060000 366.720000 9.820000 371.080000 ;
      RECT 7.060000 365.640000 9.655000 366.720000 ;
      RECT 7.060000 361.280000 9.820000 365.640000 ;
      RECT 7.060000 360.200000 9.655000 361.280000 ;
      RECT 7.060000 355.840000 9.820000 360.200000 ;
      RECT 7.060000 354.760000 9.655000 355.840000 ;
      RECT 7.060000 350.400000 9.820000 354.760000 ;
      RECT 7.060000 349.320000 9.655000 350.400000 ;
      RECT 7.060000 344.960000 9.820000 349.320000 ;
      RECT 7.060000 343.880000 9.655000 344.960000 ;
      RECT 7.060000 339.520000 9.820000 343.880000 ;
      RECT 7.060000 338.440000 9.655000 339.520000 ;
      RECT 7.060000 334.080000 9.820000 338.440000 ;
      RECT 7.060000 333.000000 9.655000 334.080000 ;
      RECT 7.060000 328.640000 9.820000 333.000000 ;
      RECT 7.060000 327.560000 9.655000 328.640000 ;
      RECT 7.060000 323.200000 9.820000 327.560000 ;
      RECT 7.060000 322.120000 9.655000 323.200000 ;
      RECT 7.060000 317.760000 9.820000 322.120000 ;
      RECT 7.060000 316.680000 9.655000 317.760000 ;
      RECT 7.060000 312.320000 9.820000 316.680000 ;
      RECT 7.060000 311.240000 9.655000 312.320000 ;
      RECT 7.060000 306.880000 9.820000 311.240000 ;
      RECT 7.060000 305.800000 9.655000 306.880000 ;
      RECT 7.060000 301.440000 9.820000 305.800000 ;
      RECT 7.060000 300.360000 9.655000 301.440000 ;
      RECT 7.060000 296.000000 9.820000 300.360000 ;
      RECT 7.060000 294.920000 9.655000 296.000000 ;
      RECT 7.060000 290.560000 9.820000 294.920000 ;
      RECT 7.060000 289.480000 9.655000 290.560000 ;
      RECT 7.060000 285.120000 9.820000 289.480000 ;
      RECT 7.060000 284.040000 9.655000 285.120000 ;
      RECT 7.060000 279.680000 9.820000 284.040000 ;
      RECT 7.060000 278.600000 9.655000 279.680000 ;
      RECT 7.060000 274.240000 9.820000 278.600000 ;
      RECT 7.060000 273.160000 9.655000 274.240000 ;
      RECT 7.060000 268.800000 9.820000 273.160000 ;
      RECT 7.060000 267.720000 9.655000 268.800000 ;
      RECT 7.060000 263.360000 9.820000 267.720000 ;
      RECT 7.060000 262.280000 9.655000 263.360000 ;
      RECT 7.060000 257.920000 9.820000 262.280000 ;
      RECT 7.060000 256.840000 9.655000 257.920000 ;
      RECT 7.060000 252.480000 9.820000 256.840000 ;
      RECT 7.060000 251.400000 9.655000 252.480000 ;
      RECT 7.060000 247.040000 9.820000 251.400000 ;
      RECT 7.060000 245.960000 9.655000 247.040000 ;
      RECT 7.060000 241.600000 9.820000 245.960000 ;
      RECT 7.060000 240.520000 9.655000 241.600000 ;
      RECT 7.060000 236.160000 9.820000 240.520000 ;
      RECT 7.060000 235.080000 9.655000 236.160000 ;
      RECT 7.060000 230.720000 9.820000 235.080000 ;
      RECT 7.060000 229.640000 9.655000 230.720000 ;
      RECT 7.060000 225.280000 9.820000 229.640000 ;
      RECT 7.060000 224.200000 9.655000 225.280000 ;
      RECT 7.060000 219.840000 9.820000 224.200000 ;
      RECT 7.060000 218.760000 9.655000 219.840000 ;
      RECT 7.060000 214.400000 9.820000 218.760000 ;
      RECT 7.060000 213.320000 9.655000 214.400000 ;
      RECT 7.060000 208.960000 9.820000 213.320000 ;
      RECT 7.060000 207.880000 9.655000 208.960000 ;
      RECT 7.060000 203.520000 9.820000 207.880000 ;
      RECT 7.060000 202.440000 9.655000 203.520000 ;
      RECT 7.060000 198.080000 9.820000 202.440000 ;
      RECT 7.060000 197.000000 9.655000 198.080000 ;
      RECT 7.060000 192.640000 9.820000 197.000000 ;
      RECT 7.060000 191.560000 9.655000 192.640000 ;
      RECT 7.060000 187.200000 9.820000 191.560000 ;
      RECT 7.060000 186.120000 9.655000 187.200000 ;
      RECT 7.060000 181.760000 9.820000 186.120000 ;
      RECT 7.060000 180.680000 9.655000 181.760000 ;
      RECT 7.060000 176.320000 9.820000 180.680000 ;
      RECT 7.060000 175.240000 9.655000 176.320000 ;
      RECT 7.060000 170.880000 9.820000 175.240000 ;
      RECT 7.060000 169.800000 9.655000 170.880000 ;
      RECT 7.060000 165.440000 9.820000 169.800000 ;
      RECT 7.060000 164.360000 9.655000 165.440000 ;
      RECT 7.060000 160.000000 9.820000 164.360000 ;
      RECT 7.060000 158.920000 9.655000 160.000000 ;
      RECT 7.060000 154.560000 9.820000 158.920000 ;
      RECT 7.060000 153.480000 9.655000 154.560000 ;
      RECT 7.060000 149.120000 9.820000 153.480000 ;
      RECT 7.060000 148.040000 9.655000 149.120000 ;
      RECT 7.060000 143.680000 9.820000 148.040000 ;
      RECT 7.060000 142.600000 9.655000 143.680000 ;
      RECT 7.060000 138.240000 9.820000 142.600000 ;
      RECT 7.060000 137.160000 9.655000 138.240000 ;
      RECT 7.060000 132.800000 9.820000 137.160000 ;
      RECT 7.060000 131.720000 9.655000 132.800000 ;
      RECT 7.060000 127.360000 9.820000 131.720000 ;
      RECT 7.060000 126.280000 9.655000 127.360000 ;
      RECT 7.060000 121.920000 9.820000 126.280000 ;
      RECT 7.060000 120.840000 9.655000 121.920000 ;
      RECT 7.060000 116.480000 9.820000 120.840000 ;
      RECT 7.060000 115.400000 9.655000 116.480000 ;
      RECT 7.060000 111.040000 9.820000 115.400000 ;
      RECT 7.060000 109.960000 9.655000 111.040000 ;
      RECT 7.060000 105.600000 9.820000 109.960000 ;
      RECT 7.060000 104.520000 9.655000 105.600000 ;
      RECT 7.060000 100.160000 9.820000 104.520000 ;
      RECT 7.060000 99.080000 9.655000 100.160000 ;
      RECT 7.060000 94.720000 9.820000 99.080000 ;
      RECT 7.060000 93.640000 9.655000 94.720000 ;
      RECT 7.060000 89.280000 9.820000 93.640000 ;
      RECT 7.060000 88.200000 9.655000 89.280000 ;
      RECT 7.060000 83.840000 9.820000 88.200000 ;
      RECT 7.060000 82.760000 9.655000 83.840000 ;
      RECT 7.060000 78.400000 9.820000 82.760000 ;
      RECT 7.060000 77.320000 9.655000 78.400000 ;
      RECT 7.060000 72.960000 9.820000 77.320000 ;
      RECT 7.060000 71.880000 9.655000 72.960000 ;
      RECT 7.060000 67.520000 9.820000 71.880000 ;
      RECT 7.060000 66.440000 9.655000 67.520000 ;
      RECT 7.060000 62.080000 9.820000 66.440000 ;
      RECT 7.060000 61.000000 9.655000 62.080000 ;
      RECT 7.060000 56.640000 9.820000 61.000000 ;
      RECT 7.060000 55.560000 9.655000 56.640000 ;
      RECT 7.060000 51.200000 9.820000 55.560000 ;
      RECT 7.060000 50.120000 9.655000 51.200000 ;
      RECT 7.060000 45.760000 9.820000 50.120000 ;
      RECT 7.060000 44.680000 9.655000 45.760000 ;
      RECT 7.060000 40.320000 9.820000 44.680000 ;
      RECT 7.060000 39.240000 9.655000 40.320000 ;
      RECT 7.060000 34.880000 9.820000 39.240000 ;
      RECT 7.060000 33.800000 9.655000 34.880000 ;
      RECT 7.060000 29.440000 9.820000 33.800000 ;
      RECT 7.060000 28.360000 9.655000 29.440000 ;
      RECT 7.060000 24.000000 9.820000 28.360000 ;
      RECT 7.060000 22.920000 9.655000 24.000000 ;
      RECT 7.060000 18.560000 9.820000 22.920000 ;
      RECT 7.060000 17.480000 9.655000 18.560000 ;
      RECT 7.060000 13.120000 9.820000 17.480000 ;
      RECT 7.060000 12.040000 9.655000 13.120000 ;
      RECT 508.620000 5.130000 543.100000 594.290000 ;
      RECT 506.620000 5.130000 506.820000 594.290000 ;
      RECT 463.620000 5.130000 504.820000 594.290000 ;
      RECT 461.620000 5.130000 461.820000 594.290000 ;
      RECT 418.620000 5.130000 459.820000 594.290000 ;
      RECT 416.620000 5.130000 416.820000 594.290000 ;
      RECT 373.620000 5.130000 414.820000 594.290000 ;
      RECT 371.620000 5.130000 371.820000 594.290000 ;
      RECT 328.620000 5.130000 369.820000 594.290000 ;
      RECT 326.620000 5.130000 326.820000 594.290000 ;
      RECT 283.620000 5.130000 324.820000 594.290000 ;
      RECT 281.620000 5.130000 281.820000 594.290000 ;
      RECT 238.620000 5.130000 279.820000 594.290000 ;
      RECT 236.620000 5.130000 236.820000 594.290000 ;
      RECT 193.620000 5.130000 234.820000 594.290000 ;
      RECT 191.620000 5.130000 191.820000 594.290000 ;
      RECT 148.620000 5.130000 189.820000 594.290000 ;
      RECT 146.620000 5.130000 146.820000 594.290000 ;
      RECT 103.620000 5.130000 144.820000 594.290000 ;
      RECT 101.620000 5.130000 101.820000 594.290000 ;
      RECT 58.620000 5.130000 99.820000 594.290000 ;
      RECT 56.620000 5.130000 56.820000 594.290000 ;
      RECT 13.620000 5.130000 54.820000 594.290000 ;
      RECT 11.620000 5.130000 11.820000 594.290000 ;
      RECT 506.620000 2.930000 543.100000 5.130000 ;
      RECT 461.620000 2.930000 504.820000 5.130000 ;
      RECT 416.620000 2.930000 459.820000 5.130000 ;
      RECT 371.620000 2.930000 414.820000 5.130000 ;
      RECT 326.620000 2.930000 369.820000 5.130000 ;
      RECT 281.620000 2.930000 324.820000 5.130000 ;
      RECT 236.620000 2.930000 279.820000 5.130000 ;
      RECT 191.620000 2.930000 234.820000 5.130000 ;
      RECT 146.620000 2.930000 189.820000 5.130000 ;
      RECT 101.620000 2.930000 144.820000 5.130000 ;
      RECT 56.620000 2.930000 99.820000 5.130000 ;
      RECT 11.620000 2.930000 54.820000 5.130000 ;
      RECT 7.060000 2.930000 9.820000 12.040000 ;
      RECT 547.100000 0.000000 550.160000 599.760000 ;
      RECT 544.900000 0.000000 545.300000 599.760000 ;
      RECT 7.060000 0.000000 543.100000 2.930000 ;
      RECT 4.860000 0.000000 5.260000 599.760000 ;
      RECT 0.000000 0.000000 3.060000 599.760000 ;
  END
END ibex_top

END LIBRARY
