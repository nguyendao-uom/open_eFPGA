##
## LEF for PtnCells ;
## created by Innovus v19.11-s128_1 on Thu Nov 25 18:55:31 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RAM_IO
  CLASS BLOCK ;
  SIZE 109.940000 BY 200.260000 ;
  FOREIGN RAM_IO 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.8162 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.973 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 8.320000 199.560000 8.700000 200.260000 ;
    END
  END N1BEG[3]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6218 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.001 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 6.940000 199.560000 7.320000 200.260000 ;
    END
  END N1BEG[2]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.746 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.1288 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 139.824 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 6.020000 199.560000 6.400000 200.260000 ;
    END
  END N1BEG[1]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3458 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.503 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 199.560000 5.480000 200.260000 ;
    END
  END N1BEG[0]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.5938 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.861 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 16.600000 199.560000 16.980000 200.260000 ;
    END
  END N2BEG[7]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.5366 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.457 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 15.680000 199.560000 16.060000 200.260000 ;
    END
  END N2BEG[6]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6057 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9205 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 14.760000 199.560000 15.140000 200.260000 ;
    END
  END N2BEG[5]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.595 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.2008 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 140.208 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 13.380000 199.560000 13.760000 200.260000 ;
    END
  END N2BEG[4]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.344 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 12.460000 199.560000 12.840000 200.260000 ;
    END
  END N2BEG[3]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.353 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.657 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 11.540000 199.560000 11.920000 200.260000 ;
    END
  END N2BEG[2]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.143 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 10.160000 199.560000 10.540000 200.260000 ;
    END
  END N2BEG[1]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2242 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.013 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 9.240000 199.560000 9.620000 200.260000 ;
    END
  END N2BEG[0]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3382 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.583 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 25.340000 199.560000 25.720000 200.260000 ;
    END
  END N2BEGb[7]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7642 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.713 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 24.420000 199.560000 24.800000 200.260000 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.145 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.617 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 23.040000 199.560000 23.420000 200.260000 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6218 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.001 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 22.120000 199.560000 22.500000 200.260000 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6046 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.915 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 21.200000 199.560000 21.580000 200.260000 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.955 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.667 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 19.820000 199.560000 20.200000 200.260000 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.955 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.667 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 18.900000 199.560000 19.280000 200.260000 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0814 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.299 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 17.980000 199.560000 18.360000 200.260000 ;
    END
  END N2BEGb[0]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5574 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.679 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 42.820000 199.560000 43.200000 200.260000 ;
    END
  END N4BEG[15]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4922 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 41.440000 199.560000 41.820000 200.260000 ;
    END
  END N4BEG[14]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.353 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.657 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 40.520000 199.560000 40.900000 200.260000 ;
    END
  END N4BEG[13]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1074 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.311 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 39.600000 199.560000 39.980000 200.260000 ;
    END
  END N4BEG[12]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.829 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.037 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 38.220000 199.560000 38.600000 200.260000 ;
    END
  END N4BEG[11]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.843 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.107 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 37.300000 199.560000 37.680000 200.260000 ;
    END
  END N4BEG[10]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3666 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 36.380000 199.560000 36.760000 200.260000 ;
    END
  END N4BEG[9]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.085 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 35.000000 199.560000 35.380000 200.260000 ;
    END
  END N4BEG[8]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9074 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.429 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 34.080000 199.560000 34.460000 200.260000 ;
    END
  END N4BEG[7]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 33.160000 199.560000 33.540000 200.260000 ;
    END
  END N4BEG[6]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 31.780000 199.560000 32.160000 200.260000 ;
    END
  END N4BEG[5]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7803 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.7935 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 30.860000 199.560000 31.240000 200.260000 ;
    END
  END N4BEG[4]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.441 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 29.940000 199.560000 30.320000 200.260000 ;
    END
  END N4BEG[3]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2102 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.943 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 28.560000 199.560000 28.940000 200.260000 ;
    END
  END N4BEG[2]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.955 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.667 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 27.640000 199.560000 28.020000 200.260000 ;
    END
  END N4BEG[1]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.645 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 26.260000 199.560000 26.640000 200.260000 ;
    END
  END N4BEG[0]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.9424 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.026 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 13.1622 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.5068 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.408 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 14.6595 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 56.6471 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.486312 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.7456 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 271.584 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 66.1763 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 335.688 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 8.320000 0.000000 8.700000 0.700000 ;
    END
  END N1END[3]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8859 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.9245 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 13.0297 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.5957 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.390645 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 13.7034 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 50.975 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.458019 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.6246 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 132.272 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 36.98 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 184.272 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.625157 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 6.940000 0.000000 7.320000 0.700000 ;
    END
  END N1END[2]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.3923 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.6625 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 39.9654 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 194.967 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.579644 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.0508 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.408 LAYER met3  ;
    ANTENNAGATEAREA 0.9915 LAYER met3  ;
    ANTENNAMAXAREACAR 42.0338 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 206.473 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.579644 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 6.020000 0.000000 6.400000 0.700000 ;
    END
  END N1END[1]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0455 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.7225 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 11.1699 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.8643 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.390645 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 11.5994 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 44.9096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.458019 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.0912 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 98.368 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 37.7715 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 195.269 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 0.000000 5.480000 0.700000 ;
    END
  END N1END[0]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.2574 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.116 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 49.0921 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 241.768 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 54.288 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 271.855 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAGATEAREA 0.3555 LAYER met4  ;
    ANTENNAMAXAREACAR 70.0709 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 365.751 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 16.600000 0.000000 16.980000 0.700000 ;
    END
  END N2MID[7]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6828 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.125 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 52.5023 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 258.252 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.545875 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.376 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 55.2803 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 275.433 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.7553 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 154.768 LAYER met4  ;
    ANTENNAGATEAREA 1.2249 LAYER met4  ;
    ANTENNAMAXAREACAR 78.7559 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 401.784 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 15.680000 0.000000 16.060000 0.700000 ;
    END
  END N2MID[6]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2994 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.251 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3555 LAYER met2  ;
    ANTENNAMAXAREACAR 54.0627 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 260.42 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.46478 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 14.760000 0.000000 15.140000 0.700000 ;
    END
  END N2MID[5]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.5285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.6695 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 105.84 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3555 LAYER met4  ;
    ANTENNAMAXAREACAR 80.1373 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 419.832 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 13.380000 0.000000 13.760000 0.700000 ;
    END
  END N2MID[4]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.1195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.0989 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 280.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2249 LAYER met4  ;
    ANTENNAMAXAREACAR 61.6158 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 308.325 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 12.460000 0.000000 12.840000 0.700000 ;
    END
  END N2MID[3]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.7251 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 277.744 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2249 LAYER met4  ;
    ANTENNAMAXAREACAR 83.8356 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 435.1 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 11.540000 0.000000 11.920000 0.700000 ;
    END
  END N2MID[2]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0591 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.1345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.1189 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 221.648 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2249 LAYER met4  ;
    ANTENNAMAXAREACAR 61.7949 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 321.28 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.999007 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 10.160000 0.000000 10.540000 0.700000 ;
    END
  END N2MID[1]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7214 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.253 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3555 LAYER met2  ;
    ANTENNAMAXAREACAR 52.1485 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 251.457 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 9.240000 0.000000 9.620000 0.700000 ;
    END
  END N2MID[0]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8085 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.7635 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 17.0186 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 66.3216 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 19.0499 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 78.2287 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.7198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.976 LAYER met4  ;
    ANTENNAGATEAREA 0.5937 LAYER met4  ;
    ANTENNAMAXAREACAR 44.6715 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 228.791 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 25.340000 0.000000 25.720000 0.700000 ;
    END
  END N2END[7]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2855 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 9.06395 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.7067 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 10.3016 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 32.381 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.5866 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 286.736 LAYER met4  ;
    ANTENNAGATEAREA 0.5937 LAYER met4  ;
    ANTENNAMAXAREACAR 100.56 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 525.09 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 24.420000 0.000000 24.800000 0.700000 ;
    END
  END N2END[6]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3171 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2965 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 7.72211 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.7785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.536 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 15.516 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 61.4194 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.9188 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 266.704 LAYER met4  ;
    ANTENNAGATEAREA 0.5937 LAYER met4  ;
    ANTENNAMAXAREACAR 102.409 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 536.843 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 23.040000 0.000000 23.420000 0.700000 ;
    END
  END N2END[5]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.8934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.005 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 30.5194 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 144.74 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 22.120000 0.000000 22.500000 0.700000 ;
    END
  END N2END[4]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3215 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 10.2151 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.3039 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 13.9924 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 53.5231 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.7098 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 244.256 LAYER met4  ;
    ANTENNAGATEAREA 0.5937 LAYER met4  ;
    ANTENNAMAXAREACAR 104.334 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 548.885 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 21.200000 0.000000 21.580000 0.700000 ;
    END
  END N2END[3]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5486 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.399 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 24.5205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 103.808 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 19.820000 0.000000 20.200000 0.700000 ;
    END
  END N2END[2]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8952 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.207 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 6.26708 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 12.8353 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.552 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.744 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 23.64 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 106.564 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.2698 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 236.576 LAYER met4  ;
    ANTENNAGATEAREA 0.5937 LAYER met4  ;
    ANTENNAMAXAREACAR 98.2059 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 505.042 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 18.900000 0.000000 19.280000 0.700000 ;
    END
  END N2END[1]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1808 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.635 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 6.80929 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.7016 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.954 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.888 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 18.2057 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 77.5558 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.9004 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 112.88 LAYER met4  ;
    ANTENNAGATEAREA 0.5937 LAYER met4  ;
    ANTENNAMAXAREACAR 53.4093 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 267.685 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 17.980000 0.000000 18.360000 0.700000 ;
    END
  END N2END[0]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0118 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.898 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2436 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.5124 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 132.144 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 50.9465 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 254.739 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.528511 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 42.820000 0.000000 43.200000 0.700000 ;
    END
  END N4END[15]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.4207 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.9955 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 66.6392 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 326.219 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 41.440000 0.000000 41.820000 0.700000 ;
    END
  END N4END[14]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5505 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.4508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 88.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 41.3922 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 200.136 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.38832 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 40.520000 0.000000 40.900000 0.700000 ;
    END
  END N4END[13]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.8325 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 165.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 61.1334 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 318.606 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 39.600000 0.000000 39.980000 0.700000 ;
    END
  END N4END[12]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0909 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2409 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.5848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.256 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 82.3583 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 428.611 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 38.220000 0.000000 38.600000 0.700000 ;
    END
  END N4END[11]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9927 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.2988 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 130.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 56.9129 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 292.315 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.732074 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 37.300000 0.000000 37.680000 0.700000 ;
    END
  END N4END[10]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7423 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.4196 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 152.512 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 60.6762 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 321.523 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.19033 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 36.380000 0.000000 36.760000 0.700000 ;
    END
  END N4END[9]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.3349 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.5665 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 69.6204 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 344.763 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 35.000000 0.000000 35.380000 0.700000 ;
    END
  END N4END[8]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.1976 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 167.328 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 105.313 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 560.716 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07583 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 34.080000 0.000000 34.460000 0.700000 ;
    END
  END N4END[7]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1273 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 100.784 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 65.1981 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 333.787 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.732074 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 33.160000 0.000000 33.540000 0.700000 ;
    END
  END N4END[6]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7305 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.4678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 285.632 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 117.252 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 608.116 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.729187 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 31.780000 0.000000 32.160000 0.700000 ;
    END
  END N4END[5]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.2138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 150.944 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 50.4311 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 255.496 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.208175 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 30.860000 0.000000 31.240000 0.700000 ;
    END
  END N4END[4]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.22 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.74 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 6.89947 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.9432 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.261 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.192 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 23.6029 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 106.102 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.1716 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 113.856 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 49.0227 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 246 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 29.940000 0.000000 30.320000 0.700000 ;
    END
  END N4END[3]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4421 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.9315 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 12.5855 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.1557 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 13.5056 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 50.1369 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.7157 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 201.616 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 48.2766 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 245.545 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 28.560000 0.000000 28.940000 0.700000 ;
    END
  END N4END[2]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.9402 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 53.872 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0707 LAYER met2  ;
    ANTENNAMAXAREACAR 16.6478 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 64.5832 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.360629 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.8788 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.824 LAYER met3  ;
    ANTENNAGATEAREA 1.2297 LAYER met3  ;
    ANTENNAMAXAREACAR 18.9888 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 77.4514 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 27.640000 0.000000 28.020000 0.700000 ;
    END
  END N4END[1]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.2122 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.803 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met2  ;
    ANTENNAMAXAREACAR 15.9324 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 60.5093 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.46478 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 26.260000 0.000000 26.640000 0.700000 ;
    END
  END N4END[0]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 7.29262 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 32.2036 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 80.720000 0.700000 81.100000 ;
    END
  END E1END[3]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 11.0158 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 51.9593 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 79.500000 0.700000 79.880000 ;
    END
  END E1END[2]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1089 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.056 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 15.6889 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 68.4048 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 77.670000 0.700000 78.050000 ;
    END
  END E1END[1]
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.368 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 9.23104 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 45.1501 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 76.450000 0.700000 76.830000 ;
    END
  END E1END[0]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8937 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.393 LAYER met3  ;
    ANTENNAMAXAREACAR 33.5901 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 171.695 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.783206 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 92.920000 0.700000 93.300000 ;
    END
  END E2MID[7]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.072 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 32.6735 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 164.075 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 91.090000 0.700000 91.470000 ;
    END
  END E2MID[6]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6787 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 35.0957 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 175.323 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 89.870000 0.700000 90.250000 ;
    END
  END E2MID[5]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 119.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 113.407 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 597.986 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via3  ;
    ANTENNADIFFAREA 1.3041 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.2145 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 50.08 LAYER met4  ;
    ANTENNAGATEAREA 1.5171 LAYER met4  ;
    ANTENNAMAXAREACAR 119.481 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 630.996 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 88.040000 0.700000 88.420000 ;
    END
  END E2MID[4]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 7.32136 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 28.9061 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 86.820000 0.700000 87.200000 ;
    END
  END E2MID[3]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.976 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 10.0351 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 47.6743 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 84.990000 0.700000 85.370000 ;
    END
  END E2MID[2]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 8.48193 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 39.0423 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 83.770000 0.700000 84.150000 ;
    END
  END E2MID[1]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 17.2885 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 81.2629 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 81.940000 0.700000 82.320000 ;
    END
  END E2MID[0]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3192 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.648 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4095 LAYER met3  ;
    ANTENNAMAXAREACAR 43.1552 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 217.977 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 104.510000 0.700000 104.890000 ;
    END
  END E2END[7]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.368 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.426 LAYER met3  ;
    ANTENNAMAXAREACAR 93.5815 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 463.581 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.440845 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 103.290000 0.700000 103.670000 ;
    END
  END E2END[6]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1624 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.528 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 42.5664 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 218.249 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 101.460000 0.700000 101.840000 ;
    END
  END E2END[5]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.69658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.512 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 39.8133 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 205.779 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 100.240000 0.700000 100.620000 ;
    END
  END E2END[4]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 19.2585 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 92.8826 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 98.410000 0.700000 98.790000 ;
    END
  END E2END[3]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 8.62341 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 39.374 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 97.190000 0.700000 97.570000 ;
    END
  END E2END[2]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.848 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 44.9054 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 228.136 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 95.360000 0.700000 95.740000 ;
    END
  END E2END[1]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4416 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.216 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 11.3937 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 54.1455 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 94.140000 0.700000 94.520000 ;
    END
  END E2END[0]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9016 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.0004 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 140.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met4  ;
    ANTENNAMAXAREACAR 129.884 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 681.858 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.85635 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 128.300000 0.700000 128.680000 ;
    END
  END EE4END[15]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.824 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 21.1026 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 101.465 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 127.080000 0.700000 127.460000 ;
    END
  END EE4END[14]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3434 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.16 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 19.3901 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 96.169 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 125.250000 0.700000 125.630000 ;
    END
  END EE4END[13]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.8432 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.296 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 55.7157 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 294.92 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 124.030000 0.700000 124.410000 ;
    END
  END EE4END[12]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.776 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 56.9608 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 298.629 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 122.200000 0.700000 122.580000 ;
    END
  END EE4END[11]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9754 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.864 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 34.5185 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 178.878 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 120.980000 0.700000 121.360000 ;
    END
  END EE4END[10]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0032 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.816 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 8.55892 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 43.7371 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 119.150000 0.700000 119.530000 ;
    END
  END EE4END[9]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.1692 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.368 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 51.0533 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 269.075 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 117.930000 0.700000 118.310000 ;
    END
  END EE4END[8]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.1336 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 48.6599 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 260.268 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 116.710000 0.700000 117.090000 ;
    END
  END EE4END[7]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 8.87911 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 42.4131 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 114.880000 0.700000 115.260000 ;
    END
  END EE4END[6]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 26.466 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 129.516 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 113.660000 0.700000 114.040000 ;
    END
  END EE4END[5]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.7336 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.9488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.864 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 23.2556 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 120.446 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 111.830000 0.700000 112.210000 ;
    END
  END EE4END[4]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1089 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.056 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 27.5766 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 132.504 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 110.610000 0.700000 110.990000 ;
    END
  END EE4END[3]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.368 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 16.1389 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 80.2392 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 108.780000 0.700000 109.160000 ;
    END
  END EE4END[2]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0224 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3555 LAYER met3  ;
    ANTENNAMAXAREACAR 10.6299 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 46.9299 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.435788 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 107.560000 0.700000 107.940000 ;
    END
  END EE4END[1]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.904 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 19.0707 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 94.0235 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 105.730000 0.700000 106.110000 ;
    END
  END EE4END[0]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 16.8115 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 78.662 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 145.990000 0.700000 146.370000 ;
    END
  END E6END[11]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.336 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 13.3308 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 67.5822 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 144.770000 0.700000 145.150000 ;
    END
  END E6END[10]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 14.8622 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 72.8873 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 143.550000 0.700000 143.930000 ;
    END
  END E6END[9]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.104 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 24.296 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 109.254 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 141.720000 0.700000 142.100000 ;
    END
  END E6END[8]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.368 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 23.9976 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 112.032 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 140.500000 0.700000 140.880000 ;
    END
  END E6END[7]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.4922 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 120.424 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.552 LAYER met3  ;
    ANTENNAMAXAREACAR 66.4251 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 330.373 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.822496 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 138.670000 0.700000 139.050000 ;
    END
  END E6END[6]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4095 LAYER met3  ;
    ANTENNAMAXAREACAR 17.4574 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 85.8965 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.359258 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 137.450000 0.700000 137.830000 ;
    END
  END E6END[5]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.7994 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 70.9843 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 369.347 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 135.620000 0.700000 136.000000 ;
    END
  END E6END[4]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7254 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.344 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.285 LAYER met3  ;
    ANTENNAMAXAREACAR 41.7522 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 201.528 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.726859 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 134.400000 0.700000 134.780000 ;
    END
  END E6END[3]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9054 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.304 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.372 LAYER met3  ;
    ANTENNAMAXAREACAR 38.0654 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 186.887 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.454475 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 132.570000 0.700000 132.950000 ;
    END
  END E6END[2]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.2324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.848 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 59.3191 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 310.534 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.986768 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.6718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 62.72 LAYER met4  ;
    ANTENNAGATEAREA 0.3555 LAYER met4  ;
    ANTENNAMAXAREACAR 92.1512 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 486.962 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.986768 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 131.350000 0.700000 131.730000 ;
    END
  END E6END[1]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9582 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.856 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.285 LAYER met3  ;
    ANTENNAMAXAREACAR 54.8913 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 269.295 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.21834 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.6504 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.88 LAYER met4  ;
    ANTENNAGATEAREA 0.8787 LAYER met4  ;
    ANTENNAMAXAREACAR 59.0456 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 293.057 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.21834 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 130.130000 0.700000 130.510000 ;
    END
  END E6END[0]
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.907 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 46.960000 0.000000 47.340000 0.700000 ;
    END
  END S1BEG[3]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.656 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 46.040000 0.000000 46.420000 0.700000 ;
    END
  END S1BEG[2]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.574 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.3968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 135.92 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 44.660000 0.000000 45.040000 0.700000 ;
    END
  END S1BEG[1]
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.8348 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 122.256 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 43.740000 0.000000 44.120000 0.700000 ;
    END
  END S1BEG[0]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.7902 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 53.725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 64.440000 0.000000 64.820000 0.700000 ;
    END
  END S2BEG[7]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.991 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 63.060000 0.000000 63.440000 0.700000 ;
    END
  END S2BEG[6]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4102 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 62.140000 0.000000 62.520000 0.700000 ;
    END
  END S2BEG[5]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.746 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.2268 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 161.68 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 61.220000 0.000000 61.600000 0.700000 ;
    END
  END S2BEG[4]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.353 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.657 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 59.840000 0.000000 60.220000 0.700000 ;
    END
  END S2BEG[3]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8475 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 58.920000 0.000000 59.300000 0.700000 ;
    END
  END S2BEG[2]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3194 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.489 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 58.000000 0.000000 58.380000 0.700000 ;
    END
  END S2BEG[1]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9317 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.919 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.0548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 134.096 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 56.620000 0.000000 57.000000 0.700000 ;
    END
  END S2BEG[0]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6694 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.239 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 55.700000 0.000000 56.080000 0.700000 ;
    END
  END S2BEGb[7]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0674 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.229 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 54.320000 0.000000 54.700000 0.700000 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.907 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 53.400000 0.000000 53.780000 0.700000 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.753 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.657 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 52.480000 0.000000 52.860000 0.700000 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.373 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 51.100000 0.000000 51.480000 0.700000 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.74 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.582 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 50.180000 0.000000 50.560000 0.700000 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0602 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.075 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 49.260000 0.000000 49.640000 0.700000 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3838 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.811 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 47.880000 0.000000 48.260000 0.700000 ;
    END
  END S2BEGb[0]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.774 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 81.460000 0.000000 81.840000 0.700000 ;
    END
  END S4BEG[15]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.585 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 80.540000 0.000000 80.920000 0.700000 ;
    END
  END S4BEG[14]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0985 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3845 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 79.620000 0.000000 80.000000 0.700000 ;
    END
  END S4BEG[13]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3838 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.811 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 78.240000 0.000000 78.620000 0.700000 ;
    END
  END S4BEG[12]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9978 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.763 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 77.320000 0.000000 77.700000 0.700000 ;
    END
  END S4BEG[11]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.315 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.349 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 75.940000 0.000000 76.320000 0.700000 ;
    END
  END S4BEG[10]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9382 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.583 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 75.020000 0.000000 75.400000 0.700000 ;
    END
  END S4BEG[9]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.347 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 74.100000 0.000000 74.480000 0.700000 ;
    END
  END S4BEG[8]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 72.720000 0.000000 73.100000 0.700000 ;
    END
  END S4BEG[7]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 71.800000 0.000000 72.180000 0.700000 ;
    END
  END S4BEG[6]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4882 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.215 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 70.880000 0.000000 71.260000 0.700000 ;
    END
  END S4BEG[5]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9543 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6635 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 69.500000 0.000000 69.880000 0.700000 ;
    END
  END S4BEG[4]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.347 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 68.580000 0.000000 68.960000 0.700000 ;
    END
  END S4BEG[3]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4102 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 67.660000 0.000000 68.040000 0.700000 ;
    END
  END S4BEG[2]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5504 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.644 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 66.280000 0.000000 66.660000 0.700000 ;
    END
  END S4BEG[1]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6694 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.239 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 65.360000 0.000000 65.740000 0.700000 ;
    END
  END S4BEG[0]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.7832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.979 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met2  ;
    ANTENNAMAXAREACAR 16.102 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 73.3125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.497308 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.7495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.464 LAYER met3  ;
    ANTENNAGATEAREA 1.2297 LAYER met3  ;
    ANTENNAMAXAREACAR 16.7115 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 76.9426 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.529836 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.4456 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 173.984 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 62.1269 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 320.021 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 46.960000 199.560000 47.340000 200.260000 ;
    END
  END S1END[3]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.183 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3145 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 9.37773 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 27.6259 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.849 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.328 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 13.6312 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 51.3849 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.3626 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 216.208 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 62.0355 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 316.697 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 46.040000 199.560000 46.420000 200.260000 ;
    END
  END S1END[2]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.3475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.5376 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.808 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9915 LAYER met4  ;
    ANTENNAMAXAREACAR 35.1158 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 176.058 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.545466 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 44.660000 199.560000 45.040000 200.260000 ;
    END
  END S1END[1]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3529 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4855 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 17.3713 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 68.0849 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 17.9485 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 72.2441 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.5925 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 228.096 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 59.2626 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 306.924 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 43.740000 199.560000 44.120000 200.260000 ;
    END
  END S1END[0]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.3438 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.322 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met2  ;
    ANTENNAMAXAREACAR 10.9748 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.5485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.324949 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.772 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.584 LAYER met3  ;
    ANTENNAGATEAREA 0.6312 LAYER met3  ;
    ANTENNAMAXAREACAR 12.1978 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 44.8109 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.38832 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.4836 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 245.872 LAYER met4  ;
    ANTENNAGATEAREA 1.2249 LAYER met4  ;
    ANTENNAMAXAREACAR 74.5982 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 390.835 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 64.440000 199.560000 64.820000 200.260000 ;
    END
  END S2MID[7]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.24 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.8504 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 107.28 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3555 LAYER met4  ;
    ANTENNAMAXAREACAR 74.4629 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 396.24 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 63.060000 199.560000 63.440000 200.260000 ;
    END
  END S2MID[6]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6421 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.9215 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 25.1374 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 121.344 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 29.2799 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 145.812 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAGATEAREA 0.3555 LAYER met4  ;
    ANTENNAMAXAREACAR 57.2351 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 301.42 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 62.140000 199.560000 62.520000 200.260000 ;
    END
  END S2MID[5]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0035 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.7385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.18263 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.1878 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 179.344 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2249 LAYER met4  ;
    ANTENNAMAXAREACAR 61.1449 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 316.962 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07583 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 61.220000 199.560000 61.600000 200.260000 ;
    END
  END S2MID[4]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.5316 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.186 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3555 LAYER met2  ;
    ANTENNAMAXAREACAR 27.0967 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 131.283 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 59.840000 199.560000 60.220000 200.260000 ;
    END
  END S2MID[3]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7498 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.031 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3555 LAYER met2  ;
    ANTENNAMAXAREACAR 25.158 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 120.348 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.376081 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 58.920000 199.560000 59.300000 200.260000 ;
    END
  END S2MID[2]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3916 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.486 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3555 LAYER met2  ;
    ANTENNAMAXAREACAR 26.6174 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 128.886 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 58.000000 199.560000 58.380000 200.260000 ;
    END
  END S2MID[1]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7699 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 23.5266 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 126.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3555 LAYER met4  ;
    ANTENNAMAXAREACAR 100.342 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 529.542 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07583 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 56.620000 199.560000 57.000000 200.260000 ;
    END
  END S2MID[0]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2353 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.9075 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 11.5355 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.3329 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 12.4557 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 45.314 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.0524 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 183.024 LAYER met4  ;
    ANTENNAGATEAREA 0.5937 LAYER met4  ;
    ANTENNAMAXAREACAR 77.096 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 407.519 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 55.700000 199.560000 56.080000 200.260000 ;
    END
  END S2END[7]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.525 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 11.9319 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.1491 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 54.320000 199.560000 54.700000 200.260000 ;
    END
  END S2END[6]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.595 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.631 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 15.7394 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 59.9877 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 53.400000 199.560000 53.780000 200.260000 ;
    END
  END S2END[5]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.3655 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 12.6469 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.51 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.328502 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 13.2335 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 48.6692 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.42052 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.4598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 168.256 LAYER met4  ;
    ANTENNAGATEAREA 0.5937 LAYER met4  ;
    ANTENNAMAXAREACAR 83.2298 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 437.817 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 52.480000 199.560000 52.860000 200.260000 ;
    END
  END S2END[4]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.0088 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.71 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 13.9776 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 51.4444 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 51.100000 199.560000 51.480000 200.260000 ;
    END
  END S2END[3]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.1496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.296 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 14.5658 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.2461 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 50.180000 199.560000 50.560000 200.260000 ;
    END
  END S2END[2]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.9918 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.615 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 16.2807 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.3007 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 49.260000 199.560000 49.640000 200.260000 ;
    END
  END S2END[1]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4315 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.1109 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.72 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 10.9841 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 39.4824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.9336 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 181.92 LAYER met4  ;
    ANTENNAGATEAREA 0.5937 LAYER met4  ;
    ANTENNAMAXAREACAR 80.0047 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 419.468 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 47.880000 199.560000 48.260000 200.260000 ;
    END
  END S2END[0]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.5088 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.298 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 34.3832 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 168.135 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 81.460000 199.560000 81.840000 200.260000 ;
    END
  END S4END[15]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1893 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.1566 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 81.776 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 31.2954 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 159.965 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.38832 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 80.540000 199.560000 80.920000 200.260000 ;
    END
  END S4END[14]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.393 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 24.1817 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 117.728 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 79.620000 199.560000 80.000000 200.260000 ;
    END
  END S4END[13]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8119 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.8985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.643 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.2058 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.568 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 55.4005 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 296.015 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 78.240000 199.560000 78.620000 200.260000 ;
    END
  END S4END[12]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.384 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 22.1369 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 107.504 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 77.320000 199.560000 77.700000 200.260000 ;
    END
  END S4END[11]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0605 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.1415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.8906 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 91.024 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 35.9506 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 182.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.502824 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 75.940000 199.560000 76.320000 200.260000 ;
    END
  END S4END[10]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5654 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.699 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 29.8361 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 145.656 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 75.020000 199.560000 75.400000 200.260000 ;
    END
  END S4END[9]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.18 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 28.0173 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 136.99 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 74.100000 199.560000 74.480000 200.260000 ;
    END
  END S4END[8]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1249 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.4006 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 61.744 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 65.033 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 348.967 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 72.720000 199.560000 73.100000 200.260000 ;
    END
  END S4END[7]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5767 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.7225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.687 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.7414 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 96.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 37.7777 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 195.124 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.38832 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 71.800000 199.560000 72.180000 200.260000 ;
    END
  END S4END[6]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5923 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.5645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 26.371 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 131.043 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 70.880000 199.560000 71.260000 200.260000 ;
    END
  END S4END[5]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9684 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.596 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 33.4214 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 163.066 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 69.500000 199.560000 69.880000 200.260000 ;
    END
  END S4END[4]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.4561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.2055 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0707 LAYER met2  ;
    ANTENNAMAXAREACAR 25.3488 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 119.623 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.643648 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAGATEAREA 1.0707 LAYER met3  ;
    ANTENNAMAXAREACAR 25.7224 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 122.051 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.681007 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.2028 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 145.552 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 47.8439 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 240.415 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 68.580000 199.560000 68.960000 200.260000 ;
    END
  END S4END[3]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.7822 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 83.125 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met2  ;
    ANTENNAMAXAREACAR 22.2023 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 105.614 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.46478 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 67.660000 199.560000 68.040000 200.260000 ;
    END
  END S4END[2]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6151 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8065 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 10.2236 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.6179 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 13.0485 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 48.7578 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.1724 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 167.664 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 38.8735 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 199.74 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.565409 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 66.280000 199.560000 66.660000 200.260000 ;
    END
  END S4END[1]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.6437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.9495 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 15.3347 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 58.1735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 19.112 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 79.3927 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.7408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 175.088 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 45.7371 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 221.775 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.423899 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 65.360000 199.560000 65.740000 200.260000 ;
    END
  END S4END[0]
  PIN W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.8864 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.056 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 9.350000 0.700000 9.730000 ;
    END
  END W1BEG[3]
  PIN W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 7.520000 0.700000 7.900000 ;
    END
  END W1BEG[2]
  PIN W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.6124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.928 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 6.300000 0.700000 6.680000 ;
    END
  END W1BEG[1]
  PIN W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 5.080000 0.700000 5.460000 ;
    END
  END W1BEG[0]
  PIN W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 20.940000 0.700000 21.320000 ;
    END
  END W2BEG[7]
  PIN W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 19.720000 0.700000 20.100000 ;
    END
  END W2BEG[6]
  PIN W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 17.890000 0.700000 18.270000 ;
    END
  END W2BEG[5]
  PIN W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.264 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 16.670000 0.700000 17.050000 ;
    END
  END W2BEG[4]
  PIN W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 15.450000 0.700000 15.830000 ;
    END
  END W2BEG[3]
  PIN W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 13.620000 0.700000 14.000000 ;
    END
  END W2BEG[2]
  PIN W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 12.400000 0.700000 12.780000 ;
    END
  END W2BEG[1]
  PIN W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.1144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.272 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 10.570000 0.700000 10.950000 ;
    END
  END W2BEG[0]
  PIN W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.6784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 33.140000 0.700000 33.520000 ;
    END
  END W2BEGb[7]
  PIN W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 31.310000 0.700000 31.690000 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 30.090000 0.700000 30.470000 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 28.870000 0.700000 29.250000 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 27.040000 0.700000 27.420000 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.9064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.496 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 25.820000 0.700000 26.200000 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 23.990000 0.700000 24.370000 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 22.770000 0.700000 23.150000 ;
    END
  END W2BEGb[0]
  PIN WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.0718 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.52 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 56.930000 0.700000 57.310000 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.4724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.848 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 55.100000 0.700000 55.480000 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 53.880000 0.700000 54.260000 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.6984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.72 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 52.660000 0.700000 53.040000 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 50.830000 0.700000 51.210000 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.7484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.32 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 49.610000 0.700000 49.990000 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9394 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.4098 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 146.656 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 47.780000 0.700000 48.160000 ;
    END
  END WW4BEG[9]
  PIN WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.1844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.312 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 46.560000 0.700000 46.940000 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 44.730000 0.700000 45.110000 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2624 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.9106 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 43.510000 0.700000 43.890000 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.0444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.232 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 42.290000 0.700000 42.670000 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 40.460000 0.700000 40.840000 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 39.240000 0.700000 39.620000 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.5394 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 37.410000 0.700000 37.790000 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.3884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 36.190000 0.700000 36.570000 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2964 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.576 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 34.360000 0.700000 34.740000 ;
    END
  END WW4BEG[0]
  PIN W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.9454 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 74.620000 0.700000 75.000000 ;
    END
  END W6BEG[11]
  PIN W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.332 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.6296 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.632 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 73.400000 0.700000 73.780000 ;
    END
  END W6BEG[10]
  PIN W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8954 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.104 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 71.570000 0.700000 71.950000 ;
    END
  END W6BEG[9]
  PIN W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7532 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.816 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 70.350000 0.700000 70.730000 ;
    END
  END W6BEG[8]
  PIN W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.9388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 208.144 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 68.520000 0.700000 68.900000 ;
    END
  END W6BEG[7]
  PIN W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 67.300000 0.700000 67.680000 ;
    END
  END W6BEG[6]
  PIN W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.0772 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.544 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 66.080000 0.700000 66.460000 ;
    END
  END W6BEG[5]
  PIN W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.6304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.024 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 64.250000 0.700000 64.630000 ;
    END
  END W6BEG[4]
  PIN W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.5956 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.9842 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 124.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 63.030000 0.700000 63.410000 ;
    END
  END W6BEG[3]
  PIN W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4766 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.2436 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.24 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 61.200000 0.700000 61.580000 ;
    END
  END W6BEG[2]
  PIN W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.8874 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.728 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 59.980000 0.700000 60.360000 ;
    END
  END W6BEG[1]
  PIN W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0976 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.5238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.264 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 58.150000 0.700000 58.530000 ;
    END
  END W6BEG[0]
  PIN RAM2FAB_D0_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.5154 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.2572 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 36.1808 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 199.54 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 33.750000 109.940000 34.130000 ;
    END
  END RAM2FAB_D0_I0
  PIN RAM2FAB_D0_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 26.2512 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 128.892 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 36.190000 109.940000 36.570000 ;
    END
  END RAM2FAB_D0_I1
  PIN RAM2FAB_D0_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.1286 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 22.5857 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 117.73 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 38.020000 109.940000 38.400000 ;
    END
  END RAM2FAB_D0_I2
  PIN RAM2FAB_D0_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.0926 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.4978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.792 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 32.4951 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 173.704 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 40.460000 109.940000 40.840000 ;
    END
  END RAM2FAB_D0_I3
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7805 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 7.9112 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.0559 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.9238 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.064 LAYER met3  ;
    ANTENNAGATEAREA 5.0427 LAYER met3  ;
    ANTENNAMAXAREACAR 8.49101 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 24.2415 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 82.840000 0.000000 83.220000 0.700000 ;
    END
  END UserCLK
  PIN RAM2FAB_D1_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.9316 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.3258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 21.0209 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 112.038 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 23.990000 109.940000 24.370000 ;
    END
  END RAM2FAB_D1_I0
  PIN RAM2FAB_D1_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.368 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.393 LAYER met3  ;
    ANTENNAMAXAREACAR 7.93893 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 37.9873 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.306107 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 26.430000 109.940000 26.810000 ;
    END
  END RAM2FAB_D1_I1
  PIN RAM2FAB_D1_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3694 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 30.2951 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 165.08 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 28.870000 109.940000 29.250000 ;
    END
  END RAM2FAB_D1_I2
  PIN RAM2FAB_D1_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.848 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 64.2921 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 320.627 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 31.310000 109.940000 31.690000 ;
    END
  END RAM2FAB_D1_I3
  PIN RAM2FAB_D2_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 10.4617 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 50.6291 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 14.230000 109.940000 14.610000 ;
    END
  END RAM2FAB_D2_I0
  PIN RAM2FAB_D2_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8556 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 52.6739 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 281.117 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 16.670000 109.940000 17.050000 ;
    END
  END RAM2FAB_D2_I1
  PIN RAM2FAB_D2_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1089 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.056 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.393 LAYER met3  ;
    ANTENNAMAXAREACAR 16.3384 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 75.1972 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.477863 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 19.110000 109.940000 19.490000 ;
    END
  END RAM2FAB_D2_I2
  PIN RAM2FAB_D2_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7996 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.6218 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 41.12 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 46.4725 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 248.408 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 21.550000 109.940000 21.930000 ;
    END
  END RAM2FAB_D2_I3
  PIN RAM2FAB_D3_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 11.9298 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 56.615 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 5.080000 109.940000 5.460000 ;
    END
  END RAM2FAB_D3_I0
  PIN RAM2FAB_D3_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4856 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.9826 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.848 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 42.0364 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 219.272 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 6.910000 109.940000 7.290000 ;
    END
  END RAM2FAB_D3_I1
  PIN RAM2FAB_D3_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 10.3293 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 49.1315 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 9.350000 109.940000 9.730000 ;
    END
  END RAM2FAB_D3_I2
  PIN RAM2FAB_D3_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.072 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 29.0969 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 145.639 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 11.790000 109.940000 12.170000 ;
    END
  END RAM2FAB_D3_I3
  PIN FAB2RAM_D0_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.4924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.288 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 110.000000 109.940000 110.380000 ;
    END
  END FAB2RAM_D0_O0
  PIN FAB2RAM_D0_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.3204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.704 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 112.440000 109.940000 112.820000 ;
    END
  END FAB2RAM_D0_O1
  PIN FAB2RAM_D0_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.9286 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.9488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.864 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 114.880000 109.940000 115.260000 ;
    END
  END FAB2RAM_D0_O2
  PIN FAB2RAM_D0_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 117.320000 109.940000 117.700000 ;
    END
  END FAB2RAM_D0_O3
  PIN FAB2RAM_D1_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 100.240000 109.940000 100.620000 ;
    END
  END FAB2RAM_D1_O0
  PIN FAB2RAM_D1_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.3174 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 102.680000 109.940000 103.060000 ;
    END
  END FAB2RAM_D1_O1
  PIN FAB2RAM_D1_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5754 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.064 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 105.120000 109.940000 105.500000 ;
    END
  END FAB2RAM_D1_O2
  PIN FAB2RAM_D1_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.8569 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.232 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 107.560000 109.940000 107.940000 ;
    END
  END FAB2RAM_D1_O3
  PIN FAB2RAM_D2_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 91.090000 109.940000 91.470000 ;
    END
  END FAB2RAM_D2_O0
  PIN FAB2RAM_D2_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.9514 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.736 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 93.530000 109.940000 93.910000 ;
    END
  END FAB2RAM_D2_O1
  PIN FAB2RAM_D2_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.6332 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.176 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 95.970000 109.940000 96.350000 ;
    END
  END FAB2RAM_D2_O2
  PIN FAB2RAM_D2_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.7464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.976 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 98.410000 109.940000 98.790000 ;
    END
  END FAB2RAM_D2_O3
  PIN FAB2RAM_D3_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.3794 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.352 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 81.330000 109.940000 81.710000 ;
    END
  END FAB2RAM_D3_O0
  PIN FAB2RAM_D3_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.1578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.312 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 83.770000 109.940000 84.150000 ;
    END
  END FAB2RAM_D3_O1
  PIN FAB2RAM_D3_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.0074 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.368 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 86.210000 109.940000 86.590000 ;
    END
  END FAB2RAM_D3_O2
  PIN FAB2RAM_D3_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4436 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.024 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.0398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 86.016 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 88.650000 109.940000 89.030000 ;
    END
  END FAB2RAM_D3_O3
  PIN FAB2RAM_A0_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.3314 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.096 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 71.570000 109.940000 71.950000 ;
    END
  END FAB2RAM_A0_O0
  PIN FAB2RAM_A0_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 74.010000 109.940000 74.390000 ;
    END
  END FAB2RAM_A0_O1
  PIN FAB2RAM_A0_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 76.450000 109.940000 76.830000 ;
    END
  END FAB2RAM_A0_O2
  PIN FAB2RAM_A0_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 78.890000 109.940000 79.270000 ;
    END
  END FAB2RAM_A0_O3
  PIN FAB2RAM_A1_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5754 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.064 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 62.420000 109.940000 62.800000 ;
    END
  END FAB2RAM_A1_O0
  PIN FAB2RAM_A1_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 64.860000 109.940000 65.240000 ;
    END
  END FAB2RAM_A1_O1
  PIN FAB2RAM_A1_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 67.300000 109.940000 67.680000 ;
    END
  END FAB2RAM_A1_O2
  PIN FAB2RAM_A1_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 69.130000 109.940000 69.510000 ;
    END
  END FAB2RAM_A1_O3
  PIN FAB2RAM_C_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.96 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 52.660000 109.940000 53.040000 ;
    END
  END FAB2RAM_C_O0
  PIN FAB2RAM_C_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.5404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.544 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 55.100000 109.940000 55.480000 ;
    END
  END FAB2RAM_C_O1
  PIN FAB2RAM_C_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 57.540000 109.940000 57.920000 ;
    END
  END FAB2RAM_C_O2
  PIN FAB2RAM_C_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3506 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.8638 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.744 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 59.980000 109.940000 60.360000 ;
    END
  END FAB2RAM_C_O3
  PIN Config_accessC_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 42.900000 109.940000 43.280000 ;
    END
  END Config_accessC_bit0
  PIN Config_accessC_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.7134 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 45.340000 109.940000 45.720000 ;
    END
  END Config_accessC_bit1
  PIN Config_accessC_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.7934 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.56 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 47.780000 109.940000 48.160000 ;
    END
  END Config_accessC_bit2
  PIN Config_accessC_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 50.220000 109.940000 50.600000 ;
    END
  END Config_accessC_bit3
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6484 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.232 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 82.840000 199.560000 83.220000 200.260000 ;
    END
  END UserCLKo
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6146 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 31.8807 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 172.848 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.875 LAYER met4  ;
    ANTENNAMAXAREACAR 74.9745 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 390.797 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 194.180000 0.700000 194.560000 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4937 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 48.7675 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 245.486 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.73505 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 28.9524 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 155.824 LAYER met4  ;
    ANTENNAGATEAREA 1.875 LAYER met4  ;
    ANTENNAMAXAREACAR 64.2088 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 328.592 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 192.350000 0.700000 192.730000 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8906 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 43.461 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 233.664 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.962 LAYER met4  ;
    ANTENNAMAXAREACAR 50.6697 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 261.716 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.13564 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 191.130000 0.700000 191.510000 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7974 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.69 LAYER met3  ;
    ANTENNAMAXAREACAR 39.2225 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 191.866 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.780202 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.5832 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 148.992 LAYER met4  ;
    ANTENNAGATEAREA 1.962 LAYER met4  ;
    ANTENNAMAXAREACAR 59.642 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 305.506 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.842138 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 189.300000 0.700000 189.680000 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 143.936 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.4685 LAYER met3  ;
    ANTENNAMAXAREACAR 63.6989 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 319.5 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.591135 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.9016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 80.416 LAYER met4  ;
    ANTENNAGATEAREA 1.9455 LAYER met4  ;
    ANTENNAMAXAREACAR 71.3585 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 360.834 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 188.080000 0.700000 188.460000 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8714 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.776 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 32.3862 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 164.025 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.2195 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 44.9175 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 242.368 LAYER met4  ;
    ANTENNAGATEAREA 1.908 LAYER met4  ;
    ANTENNAMAXAREACAR 65.0417 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 343.719 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 186.250000 0.700000 186.630000 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0846 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 57.0204 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 307.872 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9455 LAYER met4  ;
    ANTENNAMAXAREACAR 99.3777 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 515.846 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 185.030000 0.700000 185.410000 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.7556 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 55.9476 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 300.72 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9455 LAYER met4  ;
    ANTENNAMAXAREACAR 83.8122 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 440.091 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 183.200000 0.700000 183.580000 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.461 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.1213 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 156.72 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.716 LAYER met4  ;
    ANTENNAMAXAREACAR 89.1777 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 446.363 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 181.980000 0.700000 182.360000 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.5286 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.4093 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 94.256 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7865 LAYER met4  ;
    ANTENNAMAXAREACAR 52.1481 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 274.638 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 180.760000 0.700000 181.140000 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.1754 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.762 LAYER met3  ;
    ANTENNAMAXAREACAR 36.8869 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 184.63 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.62226 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 31.9446 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 171.312 LAYER met4  ;
    ANTENNAGATEAREA 1.716 LAYER met4  ;
    ANTENNAMAXAREACAR 71.0694 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 368.65 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.2195 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 178.930000 0.700000 179.310000 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.2859 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.84 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met3  ;
    ANTENNAMAXAREACAR 42.8079 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 220.242 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.700629 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 52.4106 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 282.336 LAYER met4  ;
    ANTENNAGATEAREA 1.803 LAYER met4  ;
    ANTENNAMAXAREACAR 96.9506 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 509.728 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 177.710000 0.700000 178.090000 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.9525 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.762 LAYER met3  ;
    ANTENNAMAXAREACAR 63.2608 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 320.057 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.07984 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.9912 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 55.168 LAYER met4  ;
    ANTENNAGATEAREA 1.716 LAYER met4  ;
    ANTENNAMAXAREACAR 69.0832 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 352.206 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 175.880000 0.700000 176.260000 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.9047 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 150.68 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.69 LAYER met3  ;
    ANTENNAMAXAREACAR 67.9359 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 347.459 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.47695 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 25.0269 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 135.344 LAYER met4  ;
    ANTENNAGATEAREA 1.803 LAYER met4  ;
    ANTENNAMAXAREACAR 81.8166 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 422.525 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47695 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 174.660000 0.700000 175.040000 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.7182 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.372 LAYER met3  ;
    ANTENNAMAXAREACAR 45.3692 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 235.26 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.68237 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.084 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 34.8 LAYER met4  ;
    ANTENNAGATEAREA 1.803 LAYER met4  ;
    ANTENNAMAXAREACAR 52.5334 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 266.842 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 172.830000 0.700000 173.210000 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4986 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.984 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.3016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 60.736 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2212 LAYER met4  ;
    ANTENNAMAXAREACAR 54.4077 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 286.517 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 171.610000 0.700000 171.990000 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.8923 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 117.664 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met3  ;
    ANTENNAMAXAREACAR 52.0619 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 267.218 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.636689 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.8634 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 102.016 LAYER met4  ;
    ANTENNAGATEAREA 1.7865 LAYER met4  ;
    ANTENNAMAXAREACAR 62.6207 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 324.321 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.80021 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 169.780000 0.700000 170.160000 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 46.8879 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 252.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7865 LAYER met4  ;
    ANTENNAMAXAREACAR 62.6845 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 319.336 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 168.560000 0.700000 168.940000 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5597 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.904 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met3  ;
    ANTENNAMAXAREACAR 33.4136 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 163.721 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.13564 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 38.9151 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 209.424 LAYER met4  ;
    ANTENNAGATEAREA 1.7865 LAYER met4  ;
    ANTENNAMAXAREACAR 55.1965 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 280.947 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.13564 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 167.340000 0.700000 167.720000 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5533 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.888 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.921 LAYER met3  ;
    ANTENNAMAXAREACAR 36.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 179.107 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.768828 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 28.8306 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 157.056 LAYER met4  ;
    ANTENNAGATEAREA 1.716 LAYER met4  ;
    ANTENNAMAXAREACAR 58.9551 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 305.754 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 165.510000 0.700000 165.890000 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7701 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.603 LAYER met3  ;
    ANTENNAMAXAREACAR 72.4629 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 366.506 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.3541 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.5194 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 62.848 LAYER met4  ;
    ANTENNAGATEAREA 1.716 LAYER met4  ;
    ANTENNAMAXAREACAR 79.1758 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 403.13 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.3541 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 164.290000 0.700000 164.670000 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8394 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.752 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 54.1833 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 268.524 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.53889 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.1784 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 122.048 LAYER met4  ;
    ANTENNAGATEAREA 1.716 LAYER met4  ;
    ANTENNAMAXAREACAR 67.1078 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 339.647 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.53889 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 162.460000 0.700000 162.840000 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.8691 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.376 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5607 LAYER met3  ;
    ANTENNAMAXAREACAR 38.1039 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 184.114 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.29277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.3876 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.008 LAYER met4  ;
    ANTENNAGATEAREA 2.1507 LAYER met4  ;
    ANTENNAMAXAREACAR 47.4285 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 241.846 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.29277 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 161.240000 0.700000 161.620000 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.3224 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.776 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3555 LAYER met3  ;
    ANTENNAMAXAREACAR 53.8924 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 274.674 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.885858 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 65.6937 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 355.536 LAYER met4  ;
    ANTENNAGATEAREA 1.7865 LAYER met4  ;
    ANTENNAMAXAREACAR 102.04 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 542.563 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.09371 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 159.410000 0.700000 159.790000 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3046 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.0672 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 289.76 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.716 LAYER met4  ;
    ANTENNAMAXAREACAR 105.072 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 549.81 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 158.190000 0.700000 158.570000 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6743 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.72 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 40.8415 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 208.167 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 34.0539 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 183.968 LAYER met4  ;
    ANTENNAGATEAREA 1.7865 LAYER met4  ;
    ANTENNAMAXAREACAR 67.9585 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 345.863 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 156.360000 0.700000 156.740000 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6408 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 57.8361 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 310.336 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7865 LAYER met4  ;
    ANTENNAMAXAREACAR 83.3586 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 426.182 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 155.140000 0.700000 155.520000 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.32468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 39.9193 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 195.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.936478 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 49.638 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 267.088 LAYER met4  ;
    ANTENNAGATEAREA 1.716 LAYER met4  ;
    ANTENNAMAXAREACAR 77.5231 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 398.398 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 153.920000 0.700000 154.300000 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.3222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.5283 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 102.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7865 LAYER met4  ;
    ANTENNAMAXAREACAR 43.2209 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 226.424 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.872265 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 152.090000 0.700000 152.470000 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4096 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.4492 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 174.464 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.803 LAYER met4  ;
    ANTENNAMAXAREACAR 103.608 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 544.137 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 150.870000 0.700000 151.250000 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.4926 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.7698 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 134.448 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.716 LAYER met4  ;
    ANTENNAMAXAREACAR 67.6755 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 358.812 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 149.040000 0.700000 149.420000 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4766 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 25.5465 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 139.536 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7865 LAYER met4  ;
    ANTENNAMAXAREACAR 75.4611 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 401.536 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.2195 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 147.820000 0.700000 148.200000 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 194.180000 109.940000 194.560000 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 191.740000 109.940000 192.120000 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.0674 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 189.300000 109.940000 189.680000 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 186.860000 109.940000 187.240000 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.3654 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.944 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 184.420000 109.940000 184.800000 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.4134 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.2 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 181.980000 109.940000 182.360000 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 179.540000 109.940000 179.920000 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 177.100000 109.940000 177.480000 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 174.660000 109.940000 175.040000 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 172.220000 109.940000 172.600000 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.1264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.336 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 169.780000 109.940000 170.160000 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.9734 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.52 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 167.340000 109.940000 167.720000 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.1974 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.048 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 164.900000 109.940000 165.280000 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 162.460000 109.940000 162.840000 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 160.630000 109.940000 161.010000 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 158.190000 109.940000 158.570000 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 155.750000 109.940000 156.130000 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 153.310000 109.940000 153.690000 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.656 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 150.870000 109.940000 151.250000 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 148.430000 109.940000 148.810000 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 145.990000 109.940000 146.370000 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.9214 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.576 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 143.550000 109.940000 143.930000 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 141.110000 109.940000 141.490000 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 138.670000 109.940000 139.050000 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.1264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.336 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 136.230000 109.940000 136.610000 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 133.790000 109.940000 134.170000 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 131.350000 109.940000 131.730000 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 129.520000 109.940000 129.900000 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.4494 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 127.080000 109.940000 127.460000 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.6599 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.848 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 124.640000 109.940000 125.020000 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7666 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.7918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 31.36 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 122.200000 109.940000 122.580000 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.240000 119.760000 109.940000 120.140000 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.3794 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.789 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 64.2402 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 318.206 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 104.460000 0.000000 104.840000 0.700000 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.6508 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.028 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 70.0692 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 346.323 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 103.080000 0.000000 103.460000 0.700000 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.263 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.7498 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 127.136 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 59.6599 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 312.039 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.732074 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 102.160000 0.000000 102.540000 0.700000 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.621 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.997 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 56.5476 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 279.316 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 100.780000 0.000000 101.160000 0.700000 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.9706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 74.627 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 78.3552 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 387.753 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 99.860000 0.000000 100.240000 0.700000 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9317 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.0158 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 101.888 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 55.1603 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 283.712 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.732074 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 98.940000 0.000000 99.320000 0.700000 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.3118 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 140.8 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 70.5062 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 366.767 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.732074 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 97.560000 0.000000 97.940000 0.700000 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1014 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.281 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 21.1455 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 97.0254 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 96.640000 0.000000 97.020000 0.700000 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.4275 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 131.216 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 47.7627 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 252.825 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 95.720000 0.000000 96.100000 0.700000 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.5364 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 81.424 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.4685 LAYER met2  ;
    ANTENNAMAXAREACAR 18.379 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 85.3747 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.606289 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 94.340000 0.000000 94.720000 0.700000 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.2487 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.1785 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.431 LAYER met2  ;
    ANTENNAMAXAREACAR 18.7815 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 87.6288 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.401852 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 1.431 LAYER met3  ;
    ANTENNAMAXAREACAR 18.9597 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 88.8922 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.429804 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.3078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.112 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 23.1661 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 113.65 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.779833 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 93.420000 0.000000 93.800000 0.700000 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5344 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.511 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 23.3439 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 126.848 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 51.4137 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 269.746 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 92.500000 0.000000 92.880000 0.700000 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7785 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.2717 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 119.248 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 20.3258 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 97.8914 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 91.120000 0.000000 91.500000 0.700000 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.3355 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met2  ;
    ANTENNAMAXAREACAR 38.2443 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 184.247 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.4002 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.2 LAYER met3  ;
    ANTENNAGATEAREA 2.385 LAYER met3  ;
    ANTENNAMAXAREACAR 43.0243 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 210.327 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.624109 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.7643 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 106.816 LAYER met4  ;
    ANTENNAGATEAREA 5.214 LAYER met4  ;
    ANTENNAMAXAREACAR 46.8149 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 230.813 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.05178 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 90.200000 0.000000 90.580000 0.700000 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7181 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.2035 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 26.2597 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 124.56 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.1494 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.744 LAYER met3  ;
    ANTENNAGATEAREA 1.3887 LAYER met3  ;
    ANTENNAMAXAREACAR 29.9678 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 145.258 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.632451 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.1306 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.304 LAYER met4  ;
    ANTENNAGATEAREA 5.7192 LAYER met4  ;
    ANTENNAMAXAREACAR 38.0545 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 188.491 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.632451 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 89.280000 0.000000 89.660000 0.700000 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.6991 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.8505 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.431 LAYER met2  ;
    ANTENNAMAXAREACAR 15.2371 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 70.0517 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.492732 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAGATEAREA 1.431 LAYER met3  ;
    ANTENNAMAXAREACAR 15.5648 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 72.1258 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.520685 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.0523 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.352 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 28.0244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 136.38 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.885814 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 87.900000 0.000000 88.280000 0.700000 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.8798 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.296 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met3  ;
    ANTENNAMAXAREACAR 38.5204 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 195.313 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.842138 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.6053 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 105.968 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 42.2304 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 215.365 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 86.980000 0.000000 87.360000 0.700000 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.2162 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 84.448 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.431 LAYER met2  ;
    ANTENNAMAXAREACAR 20.7705 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 98.4064 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.690147 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.26972 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.8 LAYER met3  ;
    ANTENNAGATEAREA 2.385 LAYER met3  ;
    ANTENNAMAXAREACAR 23.3993 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 112.998 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.706918 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.0086 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 38.32 LAYER met4  ;
    ANTENNAGATEAREA 5.214 LAYER met4  ;
    ANTENNAMAXAREACAR 28.0228 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 136.474 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 86.060000 0.000000 86.440000 0.700000 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2089 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.9993 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 150.736 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 41.5932 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 204.958 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 84.680000 0.000000 85.060000 0.700000 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.5579 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 57.1865 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met2  ;
    ANTENNAMAXAREACAR 26.7008 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 127.935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.407128 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.20145 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.864 LAYER met3  ;
    ANTENNAGATEAREA 1.59 LAYER met3  ;
    ANTENNAMAXAREACAR 31.2301 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 152.378 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.566128 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.4986 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.6 LAYER met4  ;
    ANTENNAGATEAREA 5.214 LAYER met4  ;
    ANTENNAMAXAREACAR 33.6272 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 165.343 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 83.760000 0.000000 84.140000 0.700000 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.1352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.45 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 104.460000 199.560000 104.840000 200.260000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8858 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.203 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 103.080000 199.560000 103.460000 200.260000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.2256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.902 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 102.160000 199.560000 102.540000 200.260000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0282 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.915 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 100.780000 199.560000 101.160000 200.260000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9382 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.583 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.860000 199.560000 100.240000 200.260000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7326 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.555 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 98.940000 199.560000 99.320000 200.260000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0605 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.1415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.2908 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.688 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 97.560000 199.560000 97.940000 200.260000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0806 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.295 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 96.640000 199.560000 97.020000 200.260000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.3964 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.756 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 95.720000 199.560000 96.100000 200.260000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.157 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.559 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 94.340000 199.560000 94.720000 200.260000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.269 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.119 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 93.420000 199.560000 93.800000 200.260000 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7814 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.799 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 92.500000 199.560000 92.880000 200.260000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.7594 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.571 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 91.120000 199.560000 91.500000 200.260000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.0658 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.221 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 90.200000 199.560000 90.580000 200.260000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.521 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.379 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 89.280000 199.560000 89.660000 200.260000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.8542 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.045 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 87.900000 199.560000 88.280000 200.260000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0282 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.915 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 86.980000 199.560000 87.360000 200.260000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3954 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.751 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 86.060000 199.560000 86.440000 200.260000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6218 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.001 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 84.680000 199.560000 85.060000 200.260000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.129 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.537 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 83.760000 199.560000 84.140000 200.260000 ;
    END
  END FrameStrobe_O[0]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 108.740000 195.020000 109.940000 196.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 195.020000 1.200000 196.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.740000 2.850000 109.940000 4.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 1.200000 4.050000 ;
    END
    PORT
      LAYER met4 ;
        RECT 105.910000 199.060000 107.110000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 105.910000 0.000000 107.110000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 199.060000 4.030000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 0.000000 4.030000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 109.940000 4.050000 ;
        RECT 0.000000 195.020000 109.940000 196.220000 ;
        RECT 2.830000 21.180000 4.030000 21.660000 ;
        RECT 2.830000 15.740000 4.030000 16.220000 ;
        RECT 2.830000 10.300000 4.030000 10.780000 ;
        RECT 2.830000 4.860000 4.030000 5.340000 ;
        RECT 2.830000 48.380000 4.030000 48.860000 ;
        RECT 2.830000 42.940000 4.030000 43.420000 ;
        RECT 2.830000 37.500000 4.030000 37.980000 ;
        RECT 2.830000 32.060000 4.030000 32.540000 ;
        RECT 2.830000 26.620000 4.030000 27.100000 ;
        RECT 7.060000 21.180000 8.260000 21.660000 ;
        RECT 7.060000 15.740000 8.260000 16.220000 ;
        RECT 7.060000 4.860000 8.260000 5.340000 ;
        RECT 7.060000 10.300000 8.260000 10.780000 ;
        RECT 52.060000 21.180000 53.260000 21.660000 ;
        RECT 52.060000 15.740000 53.260000 16.220000 ;
        RECT 52.060000 4.860000 53.260000 5.340000 ;
        RECT 52.060000 10.300000 53.260000 10.780000 ;
        RECT 7.060000 26.620000 8.260000 27.100000 ;
        RECT 7.060000 32.060000 8.260000 32.540000 ;
        RECT 7.060000 37.500000 8.260000 37.980000 ;
        RECT 7.060000 42.940000 8.260000 43.420000 ;
        RECT 7.060000 48.380000 8.260000 48.860000 ;
        RECT 52.060000 26.620000 53.260000 27.100000 ;
        RECT 52.060000 32.060000 53.260000 32.540000 ;
        RECT 52.060000 37.500000 53.260000 37.980000 ;
        RECT 52.060000 42.940000 53.260000 43.420000 ;
        RECT 52.060000 48.380000 53.260000 48.860000 ;
        RECT 2.830000 70.140000 4.030000 70.620000 ;
        RECT 2.830000 64.700000 4.030000 65.180000 ;
        RECT 2.830000 59.260000 4.030000 59.740000 ;
        RECT 2.830000 53.820000 4.030000 54.300000 ;
        RECT 2.830000 97.340000 4.030000 97.820000 ;
        RECT 2.830000 91.900000 4.030000 92.380000 ;
        RECT 2.830000 86.460000 4.030000 86.940000 ;
        RECT 2.830000 81.020000 4.030000 81.500000 ;
        RECT 2.830000 75.580000 4.030000 76.060000 ;
        RECT 7.060000 53.820000 8.260000 54.300000 ;
        RECT 7.060000 59.260000 8.260000 59.740000 ;
        RECT 7.060000 64.700000 8.260000 65.180000 ;
        RECT 7.060000 70.140000 8.260000 70.620000 ;
        RECT 52.060000 53.820000 53.260000 54.300000 ;
        RECT 52.060000 59.260000 53.260000 59.740000 ;
        RECT 52.060000 64.700000 53.260000 65.180000 ;
        RECT 52.060000 70.140000 53.260000 70.620000 ;
        RECT 7.060000 75.580000 8.260000 76.060000 ;
        RECT 7.060000 81.020000 8.260000 81.500000 ;
        RECT 7.060000 86.460000 8.260000 86.940000 ;
        RECT 7.060000 91.900000 8.260000 92.380000 ;
        RECT 7.060000 97.340000 8.260000 97.820000 ;
        RECT 52.060000 81.020000 53.260000 81.500000 ;
        RECT 52.060000 75.580000 53.260000 76.060000 ;
        RECT 52.060000 86.460000 53.260000 86.940000 ;
        RECT 52.060000 91.900000 53.260000 92.380000 ;
        RECT 52.060000 97.340000 53.260000 97.820000 ;
        RECT 97.060000 10.300000 98.260000 10.780000 ;
        RECT 97.060000 4.860000 98.260000 5.340000 ;
        RECT 97.060000 15.740000 98.260000 16.220000 ;
        RECT 97.060000 21.180000 98.260000 21.660000 ;
        RECT 97.060000 26.620000 98.260000 27.100000 ;
        RECT 97.060000 32.060000 98.260000 32.540000 ;
        RECT 97.060000 37.500000 98.260000 37.980000 ;
        RECT 97.060000 42.940000 98.260000 43.420000 ;
        RECT 97.060000 48.380000 98.260000 48.860000 ;
        RECT 105.910000 21.180000 107.110000 21.660000 ;
        RECT 105.910000 15.740000 107.110000 16.220000 ;
        RECT 105.910000 10.300000 107.110000 10.780000 ;
        RECT 105.910000 4.860000 107.110000 5.340000 ;
        RECT 105.910000 48.380000 107.110000 48.860000 ;
        RECT 105.910000 42.940000 107.110000 43.420000 ;
        RECT 105.910000 37.500000 107.110000 37.980000 ;
        RECT 105.910000 32.060000 107.110000 32.540000 ;
        RECT 105.910000 26.620000 107.110000 27.100000 ;
        RECT 97.060000 70.140000 98.260000 70.620000 ;
        RECT 97.060000 64.700000 98.260000 65.180000 ;
        RECT 97.060000 59.260000 98.260000 59.740000 ;
        RECT 97.060000 53.820000 98.260000 54.300000 ;
        RECT 97.060000 97.340000 98.260000 97.820000 ;
        RECT 97.060000 91.900000 98.260000 92.380000 ;
        RECT 97.060000 86.460000 98.260000 86.940000 ;
        RECT 97.060000 81.020000 98.260000 81.500000 ;
        RECT 97.060000 75.580000 98.260000 76.060000 ;
        RECT 105.910000 70.140000 107.110000 70.620000 ;
        RECT 105.910000 64.700000 107.110000 65.180000 ;
        RECT 105.910000 59.260000 107.110000 59.740000 ;
        RECT 105.910000 53.820000 107.110000 54.300000 ;
        RECT 105.910000 97.340000 107.110000 97.820000 ;
        RECT 105.910000 91.900000 107.110000 92.380000 ;
        RECT 105.910000 86.460000 107.110000 86.940000 ;
        RECT 105.910000 81.020000 107.110000 81.500000 ;
        RECT 105.910000 75.580000 107.110000 76.060000 ;
        RECT 2.830000 124.540000 4.030000 125.020000 ;
        RECT 2.830000 119.100000 4.030000 119.580000 ;
        RECT 2.830000 113.660000 4.030000 114.140000 ;
        RECT 2.830000 108.220000 4.030000 108.700000 ;
        RECT 2.830000 102.780000 4.030000 103.260000 ;
        RECT 2.830000 146.300000 4.030000 146.780000 ;
        RECT 2.830000 140.860000 4.030000 141.340000 ;
        RECT 2.830000 135.420000 4.030000 135.900000 ;
        RECT 2.830000 129.980000 4.030000 130.460000 ;
        RECT 7.060000 119.100000 8.260000 119.580000 ;
        RECT 7.060000 113.660000 8.260000 114.140000 ;
        RECT 7.060000 102.780000 8.260000 103.260000 ;
        RECT 7.060000 108.220000 8.260000 108.700000 ;
        RECT 7.060000 124.540000 8.260000 125.020000 ;
        RECT 52.060000 119.100000 53.260000 119.580000 ;
        RECT 52.060000 113.660000 53.260000 114.140000 ;
        RECT 52.060000 102.780000 53.260000 103.260000 ;
        RECT 52.060000 108.220000 53.260000 108.700000 ;
        RECT 52.060000 124.540000 53.260000 125.020000 ;
        RECT 7.060000 129.980000 8.260000 130.460000 ;
        RECT 7.060000 135.420000 8.260000 135.900000 ;
        RECT 7.060000 140.860000 8.260000 141.340000 ;
        RECT 7.060000 146.300000 8.260000 146.780000 ;
        RECT 52.060000 129.980000 53.260000 130.460000 ;
        RECT 52.060000 135.420000 53.260000 135.900000 ;
        RECT 52.060000 140.860000 53.260000 141.340000 ;
        RECT 52.060000 146.300000 53.260000 146.780000 ;
        RECT 2.830000 173.500000 4.030000 173.980000 ;
        RECT 2.830000 168.060000 4.030000 168.540000 ;
        RECT 2.830000 162.620000 4.030000 163.100000 ;
        RECT 2.830000 157.180000 4.030000 157.660000 ;
        RECT 2.830000 151.740000 4.030000 152.220000 ;
        RECT 2.830000 189.820000 4.030000 190.300000 ;
        RECT 2.830000 184.380000 4.030000 184.860000 ;
        RECT 2.830000 178.940000 4.030000 179.420000 ;
        RECT 7.060000 151.740000 8.260000 152.220000 ;
        RECT 7.060000 157.180000 8.260000 157.660000 ;
        RECT 7.060000 162.620000 8.260000 163.100000 ;
        RECT 7.060000 168.060000 8.260000 168.540000 ;
        RECT 7.060000 173.500000 8.260000 173.980000 ;
        RECT 52.060000 173.500000 53.260000 173.980000 ;
        RECT 52.060000 151.740000 53.260000 152.220000 ;
        RECT 52.060000 157.180000 53.260000 157.660000 ;
        RECT 52.060000 162.620000 53.260000 163.100000 ;
        RECT 52.060000 168.060000 53.260000 168.540000 ;
        RECT 7.060000 178.940000 8.260000 179.420000 ;
        RECT 7.060000 184.380000 8.260000 184.860000 ;
        RECT 7.060000 189.820000 8.260000 190.300000 ;
        RECT 52.060000 178.940000 53.260000 179.420000 ;
        RECT 52.060000 184.380000 53.260000 184.860000 ;
        RECT 52.060000 189.820000 53.260000 190.300000 ;
        RECT 97.060000 108.220000 98.260000 108.700000 ;
        RECT 97.060000 102.780000 98.260000 103.260000 ;
        RECT 97.060000 113.660000 98.260000 114.140000 ;
        RECT 97.060000 119.100000 98.260000 119.580000 ;
        RECT 97.060000 124.540000 98.260000 125.020000 ;
        RECT 97.060000 129.980000 98.260000 130.460000 ;
        RECT 97.060000 135.420000 98.260000 135.900000 ;
        RECT 97.060000 140.860000 98.260000 141.340000 ;
        RECT 97.060000 146.300000 98.260000 146.780000 ;
        RECT 105.910000 124.540000 107.110000 125.020000 ;
        RECT 105.910000 119.100000 107.110000 119.580000 ;
        RECT 105.910000 113.660000 107.110000 114.140000 ;
        RECT 105.910000 108.220000 107.110000 108.700000 ;
        RECT 105.910000 102.780000 107.110000 103.260000 ;
        RECT 105.910000 146.300000 107.110000 146.780000 ;
        RECT 105.910000 140.860000 107.110000 141.340000 ;
        RECT 105.910000 135.420000 107.110000 135.900000 ;
        RECT 105.910000 129.980000 107.110000 130.460000 ;
        RECT 97.060000 173.500000 98.260000 173.980000 ;
        RECT 97.060000 168.060000 98.260000 168.540000 ;
        RECT 97.060000 162.620000 98.260000 163.100000 ;
        RECT 97.060000 157.180000 98.260000 157.660000 ;
        RECT 97.060000 151.740000 98.260000 152.220000 ;
        RECT 97.060000 189.820000 98.260000 190.300000 ;
        RECT 97.060000 184.380000 98.260000 184.860000 ;
        RECT 97.060000 178.940000 98.260000 179.420000 ;
        RECT 105.910000 173.500000 107.110000 173.980000 ;
        RECT 105.910000 168.060000 107.110000 168.540000 ;
        RECT 105.910000 162.620000 107.110000 163.100000 ;
        RECT 105.910000 157.180000 107.110000 157.660000 ;
        RECT 105.910000 151.740000 107.110000 152.220000 ;
        RECT 105.910000 189.820000 107.110000 190.300000 ;
        RECT 105.910000 184.380000 107.110000 184.860000 ;
        RECT 105.910000 178.940000 107.110000 179.420000 ;
      LAYER met4 ;
        RECT 97.060000 2.850000 98.260000 196.220000 ;
        RECT 52.060000 2.850000 53.260000 196.220000 ;
        RECT 7.060000 2.850000 8.260000 196.220000 ;
        RECT 105.910000 0.000000 107.110000 200.260000 ;
        RECT 2.830000 0.000000 4.030000 200.260000 ;
    END
# end of P/G power stripe data as pin

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 108.740000 196.820000 109.940000 198.020000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 196.820000 1.200000 198.020000 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.740000 1.050000 109.940000 2.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 1.200000 2.250000 ;
    END
    PORT
      LAYER met4 ;
        RECT 107.710000 199.060000 108.910000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 107.710000 0.000000 108.910000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 199.060000 2.230000 200.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 0.000000 2.230000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 109.940000 2.250000 ;
        RECT 0.000000 196.820000 109.940000 198.020000 ;
        RECT 107.710000 100.060000 108.910000 100.540000 ;
        RECT 4.895000 100.060000 6.260000 100.540000 ;
        RECT 1.030000 100.060000 2.230000 100.540000 ;
        RECT 50.060000 100.060000 51.260000 100.540000 ;
        RECT 95.060000 100.060000 96.260000 100.540000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
        RECT 4.895000 45.660000 6.260000 46.140000 ;
        RECT 4.895000 29.340000 6.260000 29.820000 ;
        RECT 4.895000 34.780000 6.260000 35.260000 ;
        RECT 4.895000 40.220000 6.260000 40.700000 ;
        RECT 1.030000 23.900000 2.230000 24.380000 ;
        RECT 1.030000 18.460000 2.230000 18.940000 ;
        RECT 1.030000 13.020000 2.230000 13.500000 ;
        RECT 1.030000 7.580000 2.230000 8.060000 ;
        RECT 1.030000 45.660000 2.230000 46.140000 ;
        RECT 1.030000 40.220000 2.230000 40.700000 ;
        RECT 1.030000 34.780000 2.230000 35.260000 ;
        RECT 1.030000 29.340000 2.230000 29.820000 ;
        RECT 50.060000 23.900000 51.260000 24.380000 ;
        RECT 50.060000 18.460000 51.260000 18.940000 ;
        RECT 50.060000 13.020000 51.260000 13.500000 ;
        RECT 50.060000 7.580000 51.260000 8.060000 ;
        RECT 50.060000 45.660000 51.260000 46.140000 ;
        RECT 50.060000 40.220000 51.260000 40.700000 ;
        RECT 50.060000 34.780000 51.260000 35.260000 ;
        RECT 50.060000 29.340000 51.260000 29.820000 ;
        RECT 4.895000 51.100000 6.260000 51.580000 ;
        RECT 4.895000 56.540000 6.260000 57.020000 ;
        RECT 4.895000 61.980000 6.260000 62.460000 ;
        RECT 4.895000 67.420000 6.260000 67.900000 ;
        RECT 4.895000 72.860000 6.260000 73.340000 ;
        RECT 4.895000 94.620000 6.260000 95.100000 ;
        RECT 4.895000 89.180000 6.260000 89.660000 ;
        RECT 4.895000 78.300000 6.260000 78.780000 ;
        RECT 4.895000 83.740000 6.260000 84.220000 ;
        RECT 1.030000 72.860000 2.230000 73.340000 ;
        RECT 1.030000 67.420000 2.230000 67.900000 ;
        RECT 1.030000 61.980000 2.230000 62.460000 ;
        RECT 1.030000 56.540000 2.230000 57.020000 ;
        RECT 1.030000 51.100000 2.230000 51.580000 ;
        RECT 1.030000 94.620000 2.230000 95.100000 ;
        RECT 1.030000 89.180000 2.230000 89.660000 ;
        RECT 1.030000 83.740000 2.230000 84.220000 ;
        RECT 1.030000 78.300000 2.230000 78.780000 ;
        RECT 50.060000 72.860000 51.260000 73.340000 ;
        RECT 50.060000 67.420000 51.260000 67.900000 ;
        RECT 50.060000 61.980000 51.260000 62.460000 ;
        RECT 50.060000 56.540000 51.260000 57.020000 ;
        RECT 50.060000 51.100000 51.260000 51.580000 ;
        RECT 50.060000 94.620000 51.260000 95.100000 ;
        RECT 50.060000 89.180000 51.260000 89.660000 ;
        RECT 50.060000 83.740000 51.260000 84.220000 ;
        RECT 50.060000 78.300000 51.260000 78.780000 ;
        RECT 95.060000 23.900000 96.260000 24.380000 ;
        RECT 95.060000 18.460000 96.260000 18.940000 ;
        RECT 95.060000 13.020000 96.260000 13.500000 ;
        RECT 95.060000 7.580000 96.260000 8.060000 ;
        RECT 95.060000 45.660000 96.260000 46.140000 ;
        RECT 95.060000 40.220000 96.260000 40.700000 ;
        RECT 95.060000 34.780000 96.260000 35.260000 ;
        RECT 95.060000 29.340000 96.260000 29.820000 ;
        RECT 107.710000 23.900000 108.910000 24.380000 ;
        RECT 107.710000 18.460000 108.910000 18.940000 ;
        RECT 107.710000 13.020000 108.910000 13.500000 ;
        RECT 107.710000 7.580000 108.910000 8.060000 ;
        RECT 107.710000 45.660000 108.910000 46.140000 ;
        RECT 107.710000 40.220000 108.910000 40.700000 ;
        RECT 107.710000 34.780000 108.910000 35.260000 ;
        RECT 107.710000 29.340000 108.910000 29.820000 ;
        RECT 95.060000 72.860000 96.260000 73.340000 ;
        RECT 95.060000 67.420000 96.260000 67.900000 ;
        RECT 95.060000 61.980000 96.260000 62.460000 ;
        RECT 95.060000 51.100000 96.260000 51.580000 ;
        RECT 95.060000 56.540000 96.260000 57.020000 ;
        RECT 95.060000 94.620000 96.260000 95.100000 ;
        RECT 95.060000 89.180000 96.260000 89.660000 ;
        RECT 95.060000 83.740000 96.260000 84.220000 ;
        RECT 95.060000 78.300000 96.260000 78.780000 ;
        RECT 107.710000 72.860000 108.910000 73.340000 ;
        RECT 107.710000 67.420000 108.910000 67.900000 ;
        RECT 107.710000 61.980000 108.910000 62.460000 ;
        RECT 107.710000 56.540000 108.910000 57.020000 ;
        RECT 107.710000 51.100000 108.910000 51.580000 ;
        RECT 107.710000 94.620000 108.910000 95.100000 ;
        RECT 107.710000 89.180000 108.910000 89.660000 ;
        RECT 107.710000 83.740000 108.910000 84.220000 ;
        RECT 107.710000 78.300000 108.910000 78.780000 ;
        RECT 4.895000 105.500000 6.260000 105.980000 ;
        RECT 4.895000 110.940000 6.260000 111.420000 ;
        RECT 4.895000 116.380000 6.260000 116.860000 ;
        RECT 4.895000 121.820000 6.260000 122.300000 ;
        RECT 4.895000 149.020000 6.260000 149.500000 ;
        RECT 4.895000 143.580000 6.260000 144.060000 ;
        RECT 4.895000 127.260000 6.260000 127.740000 ;
        RECT 4.895000 132.700000 6.260000 133.180000 ;
        RECT 4.895000 138.140000 6.260000 138.620000 ;
        RECT 1.030000 121.820000 2.230000 122.300000 ;
        RECT 1.030000 116.380000 2.230000 116.860000 ;
        RECT 1.030000 110.940000 2.230000 111.420000 ;
        RECT 1.030000 105.500000 2.230000 105.980000 ;
        RECT 1.030000 149.020000 2.230000 149.500000 ;
        RECT 1.030000 143.580000 2.230000 144.060000 ;
        RECT 1.030000 138.140000 2.230000 138.620000 ;
        RECT 1.030000 132.700000 2.230000 133.180000 ;
        RECT 1.030000 127.260000 2.230000 127.740000 ;
        RECT 50.060000 121.820000 51.260000 122.300000 ;
        RECT 50.060000 116.380000 51.260000 116.860000 ;
        RECT 50.060000 110.940000 51.260000 111.420000 ;
        RECT 50.060000 105.500000 51.260000 105.980000 ;
        RECT 50.060000 149.020000 51.260000 149.500000 ;
        RECT 50.060000 143.580000 51.260000 144.060000 ;
        RECT 50.060000 138.140000 51.260000 138.620000 ;
        RECT 50.060000 132.700000 51.260000 133.180000 ;
        RECT 50.060000 127.260000 51.260000 127.740000 ;
        RECT 4.895000 154.460000 6.260000 154.940000 ;
        RECT 4.895000 159.900000 6.260000 160.380000 ;
        RECT 4.895000 165.340000 6.260000 165.820000 ;
        RECT 4.895000 170.780000 6.260000 171.260000 ;
        RECT 4.895000 192.540000 6.260000 193.020000 ;
        RECT 4.895000 176.220000 6.260000 176.700000 ;
        RECT 4.895000 181.660000 6.260000 182.140000 ;
        RECT 4.895000 187.100000 6.260000 187.580000 ;
        RECT 1.030000 170.780000 2.230000 171.260000 ;
        RECT 1.030000 165.340000 2.230000 165.820000 ;
        RECT 1.030000 154.460000 2.230000 154.940000 ;
        RECT 1.030000 159.900000 2.230000 160.380000 ;
        RECT 1.030000 192.540000 2.230000 193.020000 ;
        RECT 1.030000 187.100000 2.230000 187.580000 ;
        RECT 1.030000 181.660000 2.230000 182.140000 ;
        RECT 1.030000 176.220000 2.230000 176.700000 ;
        RECT 50.060000 170.780000 51.260000 171.260000 ;
        RECT 50.060000 165.340000 51.260000 165.820000 ;
        RECT 50.060000 159.900000 51.260000 160.380000 ;
        RECT 50.060000 154.460000 51.260000 154.940000 ;
        RECT 50.060000 192.540000 51.260000 193.020000 ;
        RECT 50.060000 187.100000 51.260000 187.580000 ;
        RECT 50.060000 176.220000 51.260000 176.700000 ;
        RECT 50.060000 181.660000 51.260000 182.140000 ;
        RECT 95.060000 121.820000 96.260000 122.300000 ;
        RECT 95.060000 116.380000 96.260000 116.860000 ;
        RECT 95.060000 105.500000 96.260000 105.980000 ;
        RECT 95.060000 110.940000 96.260000 111.420000 ;
        RECT 95.060000 149.020000 96.260000 149.500000 ;
        RECT 95.060000 143.580000 96.260000 144.060000 ;
        RECT 95.060000 138.140000 96.260000 138.620000 ;
        RECT 95.060000 132.700000 96.260000 133.180000 ;
        RECT 95.060000 127.260000 96.260000 127.740000 ;
        RECT 107.710000 121.820000 108.910000 122.300000 ;
        RECT 107.710000 116.380000 108.910000 116.860000 ;
        RECT 107.710000 110.940000 108.910000 111.420000 ;
        RECT 107.710000 105.500000 108.910000 105.980000 ;
        RECT 107.710000 149.020000 108.910000 149.500000 ;
        RECT 107.710000 143.580000 108.910000 144.060000 ;
        RECT 107.710000 138.140000 108.910000 138.620000 ;
        RECT 107.710000 132.700000 108.910000 133.180000 ;
        RECT 107.710000 127.260000 108.910000 127.740000 ;
        RECT 95.060000 170.780000 96.260000 171.260000 ;
        RECT 95.060000 165.340000 96.260000 165.820000 ;
        RECT 95.060000 154.460000 96.260000 154.940000 ;
        RECT 95.060000 159.900000 96.260000 160.380000 ;
        RECT 95.060000 192.540000 96.260000 193.020000 ;
        RECT 95.060000 187.100000 96.260000 187.580000 ;
        RECT 95.060000 181.660000 96.260000 182.140000 ;
        RECT 95.060000 176.220000 96.260000 176.700000 ;
        RECT 107.710000 170.780000 108.910000 171.260000 ;
        RECT 107.710000 165.340000 108.910000 165.820000 ;
        RECT 107.710000 154.460000 108.910000 154.940000 ;
        RECT 107.710000 159.900000 108.910000 160.380000 ;
        RECT 107.710000 192.540000 108.910000 193.020000 ;
        RECT 107.710000 187.100000 108.910000 187.580000 ;
        RECT 107.710000 181.660000 108.910000 182.140000 ;
        RECT 107.710000 176.220000 108.910000 176.700000 ;
      LAYER met4 ;
        RECT 95.060000 1.050000 96.260000 198.020000 ;
        RECT 50.060000 1.050000 51.260000 198.020000 ;
        RECT 5.060000 1.050000 6.260000 198.020000 ;
        RECT 107.710000 0.000000 108.910000 200.260000 ;
        RECT 1.030000 0.000000 2.230000 200.260000 ;
        RECT 4.895000 100.060000 6.260000 100.540000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
        RECT 4.895000 45.660000 6.260000 46.140000 ;
        RECT 4.895000 29.340000 6.260000 29.820000 ;
        RECT 4.895000 34.780000 6.260000 35.260000 ;
        RECT 4.895000 40.220000 6.260000 40.700000 ;
        RECT 4.895000 51.100000 6.260000 51.580000 ;
        RECT 4.895000 56.540000 6.260000 57.020000 ;
        RECT 4.895000 61.980000 6.260000 62.460000 ;
        RECT 4.895000 67.420000 6.260000 67.900000 ;
        RECT 4.895000 72.860000 6.260000 73.340000 ;
        RECT 4.895000 94.620000 6.260000 95.100000 ;
        RECT 4.895000 89.180000 6.260000 89.660000 ;
        RECT 4.895000 78.300000 6.260000 78.780000 ;
        RECT 4.895000 83.740000 6.260000 84.220000 ;
        RECT 4.895000 105.500000 6.260000 105.980000 ;
        RECT 4.895000 110.940000 6.260000 111.420000 ;
        RECT 4.895000 116.380000 6.260000 116.860000 ;
        RECT 4.895000 121.820000 6.260000 122.300000 ;
        RECT 4.895000 149.020000 6.260000 149.500000 ;
        RECT 4.895000 143.580000 6.260000 144.060000 ;
        RECT 4.895000 127.260000 6.260000 127.740000 ;
        RECT 4.895000 132.700000 6.260000 133.180000 ;
        RECT 4.895000 138.140000 6.260000 138.620000 ;
        RECT 4.895000 154.460000 6.260000 154.940000 ;
        RECT 4.895000 159.900000 6.260000 160.380000 ;
        RECT 4.895000 165.340000 6.260000 165.820000 ;
        RECT 4.895000 170.780000 6.260000 171.260000 ;
        RECT 4.895000 192.540000 6.260000 193.020000 ;
        RECT 4.895000 176.220000 6.260000 176.700000 ;
        RECT 4.895000 181.660000 6.260000 182.140000 ;
        RECT 4.895000 187.100000 6.260000 187.580000 ;
    END
# end of P/G power stripe data as pin

  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 109.940000 200.260000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 109.940000 200.260000 ;
    LAYER met2 ;
      RECT 104.980000 199.420000 109.940000 200.260000 ;
      RECT 103.600000 199.420000 104.320000 200.260000 ;
      RECT 102.680000 199.420000 102.940000 200.260000 ;
      RECT 101.300000 199.420000 102.020000 200.260000 ;
      RECT 100.380000 199.420000 100.640000 200.260000 ;
      RECT 99.460000 199.420000 99.720000 200.260000 ;
      RECT 98.080000 199.420000 98.800000 200.260000 ;
      RECT 97.160000 199.420000 97.420000 200.260000 ;
      RECT 96.240000 199.420000 96.500000 200.260000 ;
      RECT 94.860000 199.420000 95.580000 200.260000 ;
      RECT 93.940000 199.420000 94.200000 200.260000 ;
      RECT 93.020000 199.420000 93.280000 200.260000 ;
      RECT 91.640000 199.420000 92.360000 200.260000 ;
      RECT 90.720000 199.420000 90.980000 200.260000 ;
      RECT 89.800000 199.420000 90.060000 200.260000 ;
      RECT 88.420000 199.420000 89.140000 200.260000 ;
      RECT 87.500000 199.420000 87.760000 200.260000 ;
      RECT 86.580000 199.420000 86.840000 200.260000 ;
      RECT 85.200000 199.420000 85.920000 200.260000 ;
      RECT 84.280000 199.420000 84.540000 200.260000 ;
      RECT 83.360000 199.420000 83.620000 200.260000 ;
      RECT 81.980000 199.420000 82.700000 200.260000 ;
      RECT 81.060000 199.420000 81.320000 200.260000 ;
      RECT 80.140000 199.420000 80.400000 200.260000 ;
      RECT 78.760000 199.420000 79.480000 200.260000 ;
      RECT 77.840000 199.420000 78.100000 200.260000 ;
      RECT 76.460000 199.420000 77.180000 200.260000 ;
      RECT 75.540000 199.420000 75.800000 200.260000 ;
      RECT 74.620000 199.420000 74.880000 200.260000 ;
      RECT 73.240000 199.420000 73.960000 200.260000 ;
      RECT 72.320000 199.420000 72.580000 200.260000 ;
      RECT 71.400000 199.420000 71.660000 200.260000 ;
      RECT 70.020000 199.420000 70.740000 200.260000 ;
      RECT 69.100000 199.420000 69.360000 200.260000 ;
      RECT 68.180000 199.420000 68.440000 200.260000 ;
      RECT 66.800000 199.420000 67.520000 200.260000 ;
      RECT 65.880000 199.420000 66.140000 200.260000 ;
      RECT 64.960000 199.420000 65.220000 200.260000 ;
      RECT 63.580000 199.420000 64.300000 200.260000 ;
      RECT 62.660000 199.420000 62.920000 200.260000 ;
      RECT 61.740000 199.420000 62.000000 200.260000 ;
      RECT 60.360000 199.420000 61.080000 200.260000 ;
      RECT 59.440000 199.420000 59.700000 200.260000 ;
      RECT 58.520000 199.420000 58.780000 200.260000 ;
      RECT 57.140000 199.420000 57.860000 200.260000 ;
      RECT 56.220000 199.420000 56.480000 200.260000 ;
      RECT 54.840000 199.420000 55.560000 200.260000 ;
      RECT 53.920000 199.420000 54.180000 200.260000 ;
      RECT 53.000000 199.420000 53.260000 200.260000 ;
      RECT 51.620000 199.420000 52.340000 200.260000 ;
      RECT 50.700000 199.420000 50.960000 200.260000 ;
      RECT 49.780000 199.420000 50.040000 200.260000 ;
      RECT 48.400000 199.420000 49.120000 200.260000 ;
      RECT 47.480000 199.420000 47.740000 200.260000 ;
      RECT 46.560000 199.420000 46.820000 200.260000 ;
      RECT 45.180000 199.420000 45.900000 200.260000 ;
      RECT 44.260000 199.420000 44.520000 200.260000 ;
      RECT 43.340000 199.420000 43.600000 200.260000 ;
      RECT 41.960000 199.420000 42.680000 200.260000 ;
      RECT 41.040000 199.420000 41.300000 200.260000 ;
      RECT 40.120000 199.420000 40.380000 200.260000 ;
      RECT 38.740000 199.420000 39.460000 200.260000 ;
      RECT 37.820000 199.420000 38.080000 200.260000 ;
      RECT 36.900000 199.420000 37.160000 200.260000 ;
      RECT 35.520000 199.420000 36.240000 200.260000 ;
      RECT 34.600000 199.420000 34.860000 200.260000 ;
      RECT 33.680000 199.420000 33.940000 200.260000 ;
      RECT 32.300000 199.420000 33.020000 200.260000 ;
      RECT 31.380000 199.420000 31.640000 200.260000 ;
      RECT 30.460000 199.420000 30.720000 200.260000 ;
      RECT 29.080000 199.420000 29.800000 200.260000 ;
      RECT 28.160000 199.420000 28.420000 200.260000 ;
      RECT 26.780000 199.420000 27.500000 200.260000 ;
      RECT 25.860000 199.420000 26.120000 200.260000 ;
      RECT 24.940000 199.420000 25.200000 200.260000 ;
      RECT 23.560000 199.420000 24.280000 200.260000 ;
      RECT 22.640000 199.420000 22.900000 200.260000 ;
      RECT 21.720000 199.420000 21.980000 200.260000 ;
      RECT 20.340000 199.420000 21.060000 200.260000 ;
      RECT 19.420000 199.420000 19.680000 200.260000 ;
      RECT 18.500000 199.420000 18.760000 200.260000 ;
      RECT 17.120000 199.420000 17.840000 200.260000 ;
      RECT 16.200000 199.420000 16.460000 200.260000 ;
      RECT 15.280000 199.420000 15.540000 200.260000 ;
      RECT 13.900000 199.420000 14.620000 200.260000 ;
      RECT 12.980000 199.420000 13.240000 200.260000 ;
      RECT 12.060000 199.420000 12.320000 200.260000 ;
      RECT 10.680000 199.420000 11.400000 200.260000 ;
      RECT 9.760000 199.420000 10.020000 200.260000 ;
      RECT 8.840000 199.420000 9.100000 200.260000 ;
      RECT 7.460000 199.420000 8.180000 200.260000 ;
      RECT 6.540000 199.420000 6.800000 200.260000 ;
      RECT 5.620000 199.420000 5.880000 200.260000 ;
      RECT 0.000000 199.420000 4.960000 200.260000 ;
      RECT 0.000000 0.840000 109.940000 199.420000 ;
      RECT 104.980000 0.000000 109.940000 0.840000 ;
      RECT 103.600000 0.000000 104.320000 0.840000 ;
      RECT 102.680000 0.000000 102.940000 0.840000 ;
      RECT 101.300000 0.000000 102.020000 0.840000 ;
      RECT 100.380000 0.000000 100.640000 0.840000 ;
      RECT 99.460000 0.000000 99.720000 0.840000 ;
      RECT 98.080000 0.000000 98.800000 0.840000 ;
      RECT 97.160000 0.000000 97.420000 0.840000 ;
      RECT 96.240000 0.000000 96.500000 0.840000 ;
      RECT 94.860000 0.000000 95.580000 0.840000 ;
      RECT 93.940000 0.000000 94.200000 0.840000 ;
      RECT 93.020000 0.000000 93.280000 0.840000 ;
      RECT 91.640000 0.000000 92.360000 0.840000 ;
      RECT 90.720000 0.000000 90.980000 0.840000 ;
      RECT 89.800000 0.000000 90.060000 0.840000 ;
      RECT 88.420000 0.000000 89.140000 0.840000 ;
      RECT 87.500000 0.000000 87.760000 0.840000 ;
      RECT 86.580000 0.000000 86.840000 0.840000 ;
      RECT 85.200000 0.000000 85.920000 0.840000 ;
      RECT 84.280000 0.000000 84.540000 0.840000 ;
      RECT 83.360000 0.000000 83.620000 0.840000 ;
      RECT 81.980000 0.000000 82.700000 0.840000 ;
      RECT 81.060000 0.000000 81.320000 0.840000 ;
      RECT 80.140000 0.000000 80.400000 0.840000 ;
      RECT 78.760000 0.000000 79.480000 0.840000 ;
      RECT 77.840000 0.000000 78.100000 0.840000 ;
      RECT 76.460000 0.000000 77.180000 0.840000 ;
      RECT 75.540000 0.000000 75.800000 0.840000 ;
      RECT 74.620000 0.000000 74.880000 0.840000 ;
      RECT 73.240000 0.000000 73.960000 0.840000 ;
      RECT 72.320000 0.000000 72.580000 0.840000 ;
      RECT 71.400000 0.000000 71.660000 0.840000 ;
      RECT 70.020000 0.000000 70.740000 0.840000 ;
      RECT 69.100000 0.000000 69.360000 0.840000 ;
      RECT 68.180000 0.000000 68.440000 0.840000 ;
      RECT 66.800000 0.000000 67.520000 0.840000 ;
      RECT 65.880000 0.000000 66.140000 0.840000 ;
      RECT 64.960000 0.000000 65.220000 0.840000 ;
      RECT 63.580000 0.000000 64.300000 0.840000 ;
      RECT 62.660000 0.000000 62.920000 0.840000 ;
      RECT 61.740000 0.000000 62.000000 0.840000 ;
      RECT 60.360000 0.000000 61.080000 0.840000 ;
      RECT 59.440000 0.000000 59.700000 0.840000 ;
      RECT 58.520000 0.000000 58.780000 0.840000 ;
      RECT 57.140000 0.000000 57.860000 0.840000 ;
      RECT 56.220000 0.000000 56.480000 0.840000 ;
      RECT 54.840000 0.000000 55.560000 0.840000 ;
      RECT 53.920000 0.000000 54.180000 0.840000 ;
      RECT 53.000000 0.000000 53.260000 0.840000 ;
      RECT 51.620000 0.000000 52.340000 0.840000 ;
      RECT 50.700000 0.000000 50.960000 0.840000 ;
      RECT 49.780000 0.000000 50.040000 0.840000 ;
      RECT 48.400000 0.000000 49.120000 0.840000 ;
      RECT 47.480000 0.000000 47.740000 0.840000 ;
      RECT 46.560000 0.000000 46.820000 0.840000 ;
      RECT 45.180000 0.000000 45.900000 0.840000 ;
      RECT 44.260000 0.000000 44.520000 0.840000 ;
      RECT 43.340000 0.000000 43.600000 0.840000 ;
      RECT 41.960000 0.000000 42.680000 0.840000 ;
      RECT 41.040000 0.000000 41.300000 0.840000 ;
      RECT 40.120000 0.000000 40.380000 0.840000 ;
      RECT 38.740000 0.000000 39.460000 0.840000 ;
      RECT 37.820000 0.000000 38.080000 0.840000 ;
      RECT 36.900000 0.000000 37.160000 0.840000 ;
      RECT 35.520000 0.000000 36.240000 0.840000 ;
      RECT 34.600000 0.000000 34.860000 0.840000 ;
      RECT 33.680000 0.000000 33.940000 0.840000 ;
      RECT 32.300000 0.000000 33.020000 0.840000 ;
      RECT 31.380000 0.000000 31.640000 0.840000 ;
      RECT 30.460000 0.000000 30.720000 0.840000 ;
      RECT 29.080000 0.000000 29.800000 0.840000 ;
      RECT 28.160000 0.000000 28.420000 0.840000 ;
      RECT 26.780000 0.000000 27.500000 0.840000 ;
      RECT 25.860000 0.000000 26.120000 0.840000 ;
      RECT 24.940000 0.000000 25.200000 0.840000 ;
      RECT 23.560000 0.000000 24.280000 0.840000 ;
      RECT 22.640000 0.000000 22.900000 0.840000 ;
      RECT 21.720000 0.000000 21.980000 0.840000 ;
      RECT 20.340000 0.000000 21.060000 0.840000 ;
      RECT 19.420000 0.000000 19.680000 0.840000 ;
      RECT 18.500000 0.000000 18.760000 0.840000 ;
      RECT 17.120000 0.000000 17.840000 0.840000 ;
      RECT 16.200000 0.000000 16.460000 0.840000 ;
      RECT 15.280000 0.000000 15.540000 0.840000 ;
      RECT 13.900000 0.000000 14.620000 0.840000 ;
      RECT 12.980000 0.000000 13.240000 0.840000 ;
      RECT 12.060000 0.000000 12.320000 0.840000 ;
      RECT 10.680000 0.000000 11.400000 0.840000 ;
      RECT 9.760000 0.000000 10.020000 0.840000 ;
      RECT 8.840000 0.000000 9.100000 0.840000 ;
      RECT 7.460000 0.000000 8.180000 0.840000 ;
      RECT 6.540000 0.000000 6.800000 0.840000 ;
      RECT 5.620000 0.000000 5.880000 0.840000 ;
      RECT 0.000000 0.000000 4.960000 0.840000 ;
    LAYER met3 ;
      RECT 0.000000 198.320000 109.940000 200.260000 ;
      RECT 1.000000 193.880000 108.940000 194.720000 ;
      RECT 0.000000 193.320000 109.940000 193.880000 ;
      RECT 0.000000 193.030000 0.730000 193.320000 ;
      RECT 109.210000 192.420000 109.940000 193.320000 ;
      RECT 96.560000 192.240000 107.410000 193.320000 ;
      RECT 51.560000 192.240000 94.760000 193.320000 ;
      RECT 6.560000 192.240000 49.760000 193.320000 ;
      RECT 2.530000 192.240000 4.595000 193.320000 ;
      RECT 1.000000 192.050000 108.940000 192.240000 ;
      RECT 0.000000 191.810000 108.940000 192.050000 ;
      RECT 1.000000 191.440000 108.940000 191.810000 ;
      RECT 1.000000 190.830000 109.940000 191.440000 ;
      RECT 0.000000 190.600000 109.940000 190.830000 ;
      RECT 107.410000 189.980000 109.940000 190.600000 ;
      RECT 0.000000 189.980000 2.530000 190.600000 ;
      RECT 107.410000 189.520000 108.940000 189.980000 ;
      RECT 98.560000 189.520000 105.610000 190.600000 ;
      RECT 53.560000 189.520000 96.760000 190.600000 ;
      RECT 8.560000 189.520000 51.760000 190.600000 ;
      RECT 4.330000 189.520000 6.760000 190.600000 ;
      RECT 1.000000 189.520000 2.530000 189.980000 ;
      RECT 1.000000 189.000000 108.940000 189.520000 ;
      RECT 0.000000 188.760000 109.940000 189.000000 ;
      RECT 1.000000 187.880000 109.940000 188.760000 ;
      RECT 109.210000 187.540000 109.940000 187.880000 ;
      RECT 0.000000 186.930000 0.730000 187.780000 ;
      RECT 96.560000 186.800000 107.410000 187.880000 ;
      RECT 51.560000 186.800000 94.760000 187.880000 ;
      RECT 6.560000 186.800000 49.760000 187.880000 ;
      RECT 2.530000 186.800000 4.595000 187.880000 ;
      RECT 1.000000 186.560000 108.940000 186.800000 ;
      RECT 1.000000 185.950000 109.940000 186.560000 ;
      RECT 0.000000 185.710000 109.940000 185.950000 ;
      RECT 1.000000 185.160000 109.940000 185.710000 ;
      RECT 107.410000 185.100000 109.940000 185.160000 ;
      RECT 1.000000 184.730000 2.530000 185.160000 ;
      RECT 107.410000 184.120000 108.940000 185.100000 ;
      RECT 107.410000 184.080000 109.940000 184.120000 ;
      RECT 98.560000 184.080000 105.610000 185.160000 ;
      RECT 53.560000 184.080000 96.760000 185.160000 ;
      RECT 8.560000 184.080000 51.760000 185.160000 ;
      RECT 4.330000 184.080000 6.760000 185.160000 ;
      RECT 0.000000 184.080000 2.530000 184.730000 ;
      RECT 0.000000 183.880000 109.940000 184.080000 ;
      RECT 1.000000 182.900000 109.940000 183.880000 ;
      RECT 0.000000 182.660000 109.940000 182.900000 ;
      RECT 1.000000 182.440000 108.940000 182.660000 ;
      RECT 0.000000 181.440000 0.730000 181.680000 ;
      RECT 109.210000 181.360000 109.940000 181.680000 ;
      RECT 96.560000 181.360000 107.410000 182.440000 ;
      RECT 51.560000 181.360000 94.760000 182.440000 ;
      RECT 6.560000 181.360000 49.760000 182.440000 ;
      RECT 2.530000 181.360000 4.595000 182.440000 ;
      RECT 1.000000 180.460000 109.940000 181.360000 ;
      RECT 0.000000 180.220000 109.940000 180.460000 ;
      RECT 0.000000 179.720000 108.940000 180.220000 ;
      RECT 0.000000 179.610000 2.530000 179.720000 ;
      RECT 107.410000 179.240000 108.940000 179.720000 ;
      RECT 107.410000 178.640000 109.940000 179.240000 ;
      RECT 98.560000 178.640000 105.610000 179.720000 ;
      RECT 53.560000 178.640000 96.760000 179.720000 ;
      RECT 8.560000 178.640000 51.760000 179.720000 ;
      RECT 4.330000 178.640000 6.760000 179.720000 ;
      RECT 1.000000 178.640000 2.530000 179.610000 ;
      RECT 1.000000 178.630000 109.940000 178.640000 ;
      RECT 0.000000 178.390000 109.940000 178.630000 ;
      RECT 1.000000 177.780000 109.940000 178.390000 ;
      RECT 1.000000 177.410000 108.940000 177.780000 ;
      RECT 0.000000 177.000000 108.940000 177.410000 ;
      RECT 0.000000 176.560000 0.730000 177.000000 ;
      RECT 109.210000 175.920000 109.940000 176.800000 ;
      RECT 96.560000 175.920000 107.410000 177.000000 ;
      RECT 51.560000 175.920000 94.760000 177.000000 ;
      RECT 6.560000 175.920000 49.760000 177.000000 ;
      RECT 2.530000 175.920000 4.595000 177.000000 ;
      RECT 1.000000 175.580000 109.940000 175.920000 ;
      RECT 0.000000 175.340000 109.940000 175.580000 ;
      RECT 1.000000 174.360000 108.940000 175.340000 ;
      RECT 0.000000 174.280000 109.940000 174.360000 ;
      RECT 0.000000 173.510000 2.530000 174.280000 ;
      RECT 107.410000 173.200000 109.940000 174.280000 ;
      RECT 98.560000 173.200000 105.610000 174.280000 ;
      RECT 53.560000 173.200000 96.760000 174.280000 ;
      RECT 8.560000 173.200000 51.760000 174.280000 ;
      RECT 4.330000 173.200000 6.760000 174.280000 ;
      RECT 1.000000 173.200000 2.530000 173.510000 ;
      RECT 1.000000 172.900000 109.940000 173.200000 ;
      RECT 1.000000 172.530000 108.940000 172.900000 ;
      RECT 0.000000 172.290000 108.940000 172.530000 ;
      RECT 1.000000 171.920000 108.940000 172.290000 ;
      RECT 1.000000 171.560000 109.940000 171.920000 ;
      RECT 109.210000 170.480000 109.940000 171.560000 ;
      RECT 96.560000 170.480000 107.410000 171.560000 ;
      RECT 51.560000 170.480000 94.760000 171.560000 ;
      RECT 6.560000 170.480000 49.760000 171.560000 ;
      RECT 2.530000 170.480000 4.595000 171.560000 ;
      RECT 0.000000 170.480000 0.730000 171.310000 ;
      RECT 0.000000 170.460000 109.940000 170.480000 ;
      RECT 1.000000 169.480000 108.940000 170.460000 ;
      RECT 0.000000 169.240000 109.940000 169.480000 ;
      RECT 1.000000 168.840000 109.940000 169.240000 ;
      RECT 1.000000 168.260000 2.530000 168.840000 ;
      RECT 107.410000 168.020000 109.940000 168.840000 ;
      RECT 0.000000 168.020000 2.530000 168.260000 ;
      RECT 107.410000 167.760000 108.940000 168.020000 ;
      RECT 98.560000 167.760000 105.610000 168.840000 ;
      RECT 53.560000 167.760000 96.760000 168.840000 ;
      RECT 8.560000 167.760000 51.760000 168.840000 ;
      RECT 4.330000 167.760000 6.760000 168.840000 ;
      RECT 1.000000 167.760000 2.530000 168.020000 ;
      RECT 1.000000 167.040000 108.940000 167.760000 ;
      RECT 0.000000 166.190000 109.940000 167.040000 ;
      RECT 1.000000 166.120000 109.940000 166.190000 ;
      RECT 109.210000 165.580000 109.940000 166.120000 ;
      RECT 96.560000 165.040000 107.410000 166.120000 ;
      RECT 51.560000 165.040000 94.760000 166.120000 ;
      RECT 6.560000 165.040000 49.760000 166.120000 ;
      RECT 2.530000 165.040000 4.595000 166.120000 ;
      RECT 0.000000 165.040000 0.730000 165.210000 ;
      RECT 0.000000 164.970000 108.940000 165.040000 ;
      RECT 1.000000 164.600000 108.940000 164.970000 ;
      RECT 1.000000 163.990000 109.940000 164.600000 ;
      RECT 0.000000 163.400000 109.940000 163.990000 ;
      RECT 107.410000 163.140000 109.940000 163.400000 ;
      RECT 0.000000 163.140000 2.530000 163.400000 ;
      RECT 107.410000 162.320000 108.940000 163.140000 ;
      RECT 98.560000 162.320000 105.610000 163.400000 ;
      RECT 53.560000 162.320000 96.760000 163.400000 ;
      RECT 8.560000 162.320000 51.760000 163.400000 ;
      RECT 4.330000 162.320000 6.760000 163.400000 ;
      RECT 1.000000 162.320000 2.530000 163.140000 ;
      RECT 1.000000 162.160000 108.940000 162.320000 ;
      RECT 0.000000 161.920000 109.940000 162.160000 ;
      RECT 1.000000 161.310000 109.940000 161.920000 ;
      RECT 1.000000 160.940000 108.940000 161.310000 ;
      RECT 0.000000 160.680000 108.940000 160.940000 ;
      RECT 0.000000 160.090000 0.730000 160.680000 ;
      RECT 109.210000 159.600000 109.940000 160.330000 ;
      RECT 96.560000 159.600000 107.410000 160.680000 ;
      RECT 51.560000 159.600000 94.760000 160.680000 ;
      RECT 6.560000 159.600000 49.760000 160.680000 ;
      RECT 2.530000 159.600000 4.595000 160.680000 ;
      RECT 1.000000 159.110000 109.940000 159.600000 ;
      RECT 0.000000 158.870000 109.940000 159.110000 ;
      RECT 1.000000 157.960000 108.940000 158.870000 ;
      RECT 107.410000 157.890000 108.940000 157.960000 ;
      RECT 1.000000 157.890000 2.530000 157.960000 ;
      RECT 0.000000 157.040000 2.530000 157.890000 ;
      RECT 107.410000 156.880000 109.940000 157.890000 ;
      RECT 98.560000 156.880000 105.610000 157.960000 ;
      RECT 53.560000 156.880000 96.760000 157.960000 ;
      RECT 8.560000 156.880000 51.760000 157.960000 ;
      RECT 4.330000 156.880000 6.760000 157.960000 ;
      RECT 1.000000 156.880000 2.530000 157.040000 ;
      RECT 1.000000 156.430000 109.940000 156.880000 ;
      RECT 1.000000 156.060000 108.940000 156.430000 ;
      RECT 0.000000 155.820000 108.940000 156.060000 ;
      RECT 1.000000 155.450000 108.940000 155.820000 ;
      RECT 1.000000 155.240000 109.940000 155.450000 ;
      RECT 0.000000 154.600000 0.730000 154.840000 ;
      RECT 109.210000 154.160000 109.940000 155.240000 ;
      RECT 96.560000 154.160000 107.410000 155.240000 ;
      RECT 51.560000 154.160000 94.760000 155.240000 ;
      RECT 6.560000 154.160000 49.760000 155.240000 ;
      RECT 2.530000 154.160000 4.595000 155.240000 ;
      RECT 1.000000 153.990000 109.940000 154.160000 ;
      RECT 1.000000 153.620000 108.940000 153.990000 ;
      RECT 0.000000 153.010000 108.940000 153.620000 ;
      RECT 0.000000 152.770000 109.940000 153.010000 ;
      RECT 1.000000 152.520000 109.940000 152.770000 ;
      RECT 1.000000 151.790000 2.530000 152.520000 ;
      RECT 107.410000 151.550000 109.940000 152.520000 ;
      RECT 0.000000 151.550000 2.530000 151.790000 ;
      RECT 107.410000 151.440000 108.940000 151.550000 ;
      RECT 98.560000 151.440000 105.610000 152.520000 ;
      RECT 53.560000 151.440000 96.760000 152.520000 ;
      RECT 8.560000 151.440000 51.760000 152.520000 ;
      RECT 4.330000 151.440000 6.760000 152.520000 ;
      RECT 1.000000 151.440000 2.530000 151.550000 ;
      RECT 1.000000 150.570000 108.940000 151.440000 ;
      RECT 0.000000 149.800000 109.940000 150.570000 ;
      RECT 0.000000 149.720000 0.730000 149.800000 ;
      RECT 109.210000 149.110000 109.940000 149.800000 ;
      RECT 96.560000 148.720000 107.410000 149.800000 ;
      RECT 51.560000 148.720000 94.760000 149.800000 ;
      RECT 6.560000 148.720000 49.760000 149.800000 ;
      RECT 2.530000 148.720000 4.595000 149.800000 ;
      RECT 0.000000 148.720000 0.730000 148.740000 ;
      RECT 0.000000 148.500000 108.940000 148.720000 ;
      RECT 1.000000 148.130000 108.940000 148.500000 ;
      RECT 1.000000 147.520000 109.940000 148.130000 ;
      RECT 0.000000 147.080000 109.940000 147.520000 ;
      RECT 107.410000 146.670000 109.940000 147.080000 ;
      RECT 0.000000 146.670000 2.530000 147.080000 ;
      RECT 107.410000 146.000000 108.940000 146.670000 ;
      RECT 98.560000 146.000000 105.610000 147.080000 ;
      RECT 53.560000 146.000000 96.760000 147.080000 ;
      RECT 8.560000 146.000000 51.760000 147.080000 ;
      RECT 4.330000 146.000000 6.760000 147.080000 ;
      RECT 1.000000 146.000000 2.530000 146.670000 ;
      RECT 1.000000 145.690000 108.940000 146.000000 ;
      RECT 0.000000 145.450000 109.940000 145.690000 ;
      RECT 1.000000 144.470000 109.940000 145.450000 ;
      RECT 0.000000 144.360000 109.940000 144.470000 ;
      RECT 109.210000 144.230000 109.940000 144.360000 ;
      RECT 0.000000 144.230000 0.730000 144.360000 ;
      RECT 96.560000 143.280000 107.410000 144.360000 ;
      RECT 51.560000 143.280000 94.760000 144.360000 ;
      RECT 6.560000 143.280000 49.760000 144.360000 ;
      RECT 2.530000 143.280000 4.595000 144.360000 ;
      RECT 1.000000 143.250000 108.940000 143.280000 ;
      RECT 0.000000 142.400000 109.940000 143.250000 ;
      RECT 1.000000 141.790000 109.940000 142.400000 ;
      RECT 1.000000 141.640000 108.940000 141.790000 ;
      RECT 1.000000 141.420000 2.530000 141.640000 ;
      RECT 0.000000 141.180000 2.530000 141.420000 ;
      RECT 107.410000 140.810000 108.940000 141.640000 ;
      RECT 107.410000 140.560000 109.940000 140.810000 ;
      RECT 98.560000 140.560000 105.610000 141.640000 ;
      RECT 53.560000 140.560000 96.760000 141.640000 ;
      RECT 8.560000 140.560000 51.760000 141.640000 ;
      RECT 4.330000 140.560000 6.760000 141.640000 ;
      RECT 1.000000 140.560000 2.530000 141.180000 ;
      RECT 1.000000 140.200000 109.940000 140.560000 ;
      RECT 0.000000 139.350000 109.940000 140.200000 ;
      RECT 1.000000 138.920000 108.940000 139.350000 ;
      RECT 0.000000 138.130000 0.730000 138.370000 ;
      RECT 109.210000 137.840000 109.940000 138.370000 ;
      RECT 96.560000 137.840000 107.410000 138.920000 ;
      RECT 51.560000 137.840000 94.760000 138.920000 ;
      RECT 6.560000 137.840000 49.760000 138.920000 ;
      RECT 2.530000 137.840000 4.595000 138.920000 ;
      RECT 1.000000 137.150000 109.940000 137.840000 ;
      RECT 0.000000 136.910000 109.940000 137.150000 ;
      RECT 0.000000 136.300000 108.940000 136.910000 ;
      RECT 1.000000 136.200000 108.940000 136.300000 ;
      RECT 107.410000 135.930000 108.940000 136.200000 ;
      RECT 1.000000 135.320000 2.530000 136.200000 ;
      RECT 107.410000 135.120000 109.940000 135.930000 ;
      RECT 98.560000 135.120000 105.610000 136.200000 ;
      RECT 53.560000 135.120000 96.760000 136.200000 ;
      RECT 8.560000 135.120000 51.760000 136.200000 ;
      RECT 4.330000 135.120000 6.760000 136.200000 ;
      RECT 0.000000 135.120000 2.530000 135.320000 ;
      RECT 0.000000 135.080000 109.940000 135.120000 ;
      RECT 1.000000 134.470000 109.940000 135.080000 ;
      RECT 1.000000 134.100000 108.940000 134.470000 ;
      RECT 0.000000 133.490000 108.940000 134.100000 ;
      RECT 0.000000 133.480000 109.940000 133.490000 ;
      RECT 0.000000 133.250000 0.730000 133.480000 ;
      RECT 109.210000 132.400000 109.940000 133.480000 ;
      RECT 96.560000 132.400000 107.410000 133.480000 ;
      RECT 51.560000 132.400000 94.760000 133.480000 ;
      RECT 6.560000 132.400000 49.760000 133.480000 ;
      RECT 2.530000 132.400000 4.595000 133.480000 ;
      RECT 1.000000 132.270000 109.940000 132.400000 ;
      RECT 0.000000 132.030000 109.940000 132.270000 ;
      RECT 1.000000 131.050000 108.940000 132.030000 ;
      RECT 0.000000 130.810000 109.940000 131.050000 ;
      RECT 1.000000 130.760000 109.940000 130.810000 ;
      RECT 107.410000 130.200000 109.940000 130.760000 ;
      RECT 1.000000 129.830000 2.530000 130.760000 ;
      RECT 107.410000 129.680000 108.940000 130.200000 ;
      RECT 98.560000 129.680000 105.610000 130.760000 ;
      RECT 53.560000 129.680000 96.760000 130.760000 ;
      RECT 8.560000 129.680000 51.760000 130.760000 ;
      RECT 4.330000 129.680000 6.760000 130.760000 ;
      RECT 0.000000 129.680000 2.530000 129.830000 ;
      RECT 0.000000 129.220000 108.940000 129.680000 ;
      RECT 0.000000 128.980000 109.940000 129.220000 ;
      RECT 1.000000 128.040000 109.940000 128.980000 ;
      RECT 109.210000 127.760000 109.940000 128.040000 ;
      RECT 0.000000 127.760000 0.730000 128.000000 ;
      RECT 96.560000 126.960000 107.410000 128.040000 ;
      RECT 51.560000 126.960000 94.760000 128.040000 ;
      RECT 6.560000 126.960000 49.760000 128.040000 ;
      RECT 2.530000 126.960000 4.595000 128.040000 ;
      RECT 1.000000 126.780000 108.940000 126.960000 ;
      RECT 0.000000 125.930000 109.940000 126.780000 ;
      RECT 1.000000 125.320000 109.940000 125.930000 ;
      RECT 1.000000 124.950000 2.530000 125.320000 ;
      RECT 0.000000 124.710000 2.530000 124.950000 ;
      RECT 107.410000 124.340000 108.940000 125.320000 ;
      RECT 107.410000 124.240000 109.940000 124.340000 ;
      RECT 98.560000 124.240000 105.610000 125.320000 ;
      RECT 53.560000 124.240000 96.760000 125.320000 ;
      RECT 8.560000 124.240000 51.760000 125.320000 ;
      RECT 4.330000 124.240000 6.760000 125.320000 ;
      RECT 1.000000 124.240000 2.530000 124.710000 ;
      RECT 1.000000 123.730000 109.940000 124.240000 ;
      RECT 0.000000 122.880000 109.940000 123.730000 ;
      RECT 1.000000 122.600000 108.940000 122.880000 ;
      RECT 0.000000 121.660000 0.730000 121.900000 ;
      RECT 109.210000 121.520000 109.940000 121.900000 ;
      RECT 96.560000 121.520000 107.410000 122.600000 ;
      RECT 51.560000 121.520000 94.760000 122.600000 ;
      RECT 6.560000 121.520000 49.760000 122.600000 ;
      RECT 2.530000 121.520000 4.595000 122.600000 ;
      RECT 1.000000 120.680000 109.940000 121.520000 ;
      RECT 0.000000 120.440000 109.940000 120.680000 ;
      RECT 0.000000 119.880000 108.940000 120.440000 ;
      RECT 0.000000 119.830000 2.530000 119.880000 ;
      RECT 107.410000 119.460000 108.940000 119.880000 ;
      RECT 1.000000 118.850000 2.530000 119.830000 ;
      RECT 107.410000 118.800000 109.940000 119.460000 ;
      RECT 98.560000 118.800000 105.610000 119.880000 ;
      RECT 53.560000 118.800000 96.760000 119.880000 ;
      RECT 8.560000 118.800000 51.760000 119.880000 ;
      RECT 4.330000 118.800000 6.760000 119.880000 ;
      RECT 0.000000 118.800000 2.530000 118.850000 ;
      RECT 0.000000 118.610000 109.940000 118.800000 ;
      RECT 1.000000 118.000000 109.940000 118.610000 ;
      RECT 1.000000 117.630000 108.940000 118.000000 ;
      RECT 0.000000 117.390000 108.940000 117.630000 ;
      RECT 1.000000 117.160000 108.940000 117.390000 ;
      RECT 109.210000 116.080000 109.940000 117.020000 ;
      RECT 96.560000 116.080000 107.410000 117.160000 ;
      RECT 51.560000 116.080000 94.760000 117.160000 ;
      RECT 6.560000 116.080000 49.760000 117.160000 ;
      RECT 2.530000 116.080000 4.595000 117.160000 ;
      RECT 0.000000 116.080000 0.730000 116.410000 ;
      RECT 0.000000 115.560000 109.940000 116.080000 ;
      RECT 1.000000 114.580000 108.940000 115.560000 ;
      RECT 0.000000 114.440000 109.940000 114.580000 ;
      RECT 0.000000 114.340000 2.530000 114.440000 ;
      RECT 107.410000 113.360000 109.940000 114.440000 ;
      RECT 98.560000 113.360000 105.610000 114.440000 ;
      RECT 53.560000 113.360000 96.760000 114.440000 ;
      RECT 8.560000 113.360000 51.760000 114.440000 ;
      RECT 4.330000 113.360000 6.760000 114.440000 ;
      RECT 1.000000 113.360000 2.530000 114.340000 ;
      RECT 0.000000 113.120000 109.940000 113.360000 ;
      RECT 0.000000 112.510000 108.940000 113.120000 ;
      RECT 1.000000 112.140000 108.940000 112.510000 ;
      RECT 1.000000 111.720000 109.940000 112.140000 ;
      RECT 0.000000 111.290000 0.730000 111.530000 ;
      RECT 109.210000 110.680000 109.940000 111.720000 ;
      RECT 96.560000 110.640000 107.410000 111.720000 ;
      RECT 51.560000 110.640000 94.760000 111.720000 ;
      RECT 6.560000 110.640000 49.760000 111.720000 ;
      RECT 2.530000 110.640000 4.595000 111.720000 ;
      RECT 1.000000 110.310000 108.940000 110.640000 ;
      RECT 0.000000 109.700000 108.940000 110.310000 ;
      RECT 0.000000 109.460000 109.940000 109.700000 ;
      RECT 1.000000 109.000000 109.940000 109.460000 ;
      RECT 1.000000 108.480000 2.530000 109.000000 ;
      RECT 107.410000 108.240000 109.940000 109.000000 ;
      RECT 0.000000 108.240000 2.530000 108.480000 ;
      RECT 107.410000 107.920000 108.940000 108.240000 ;
      RECT 98.560000 107.920000 105.610000 109.000000 ;
      RECT 53.560000 107.920000 96.760000 109.000000 ;
      RECT 8.560000 107.920000 51.760000 109.000000 ;
      RECT 4.330000 107.920000 6.760000 109.000000 ;
      RECT 1.000000 107.920000 2.530000 108.240000 ;
      RECT 1.000000 107.260000 108.940000 107.920000 ;
      RECT 0.000000 106.410000 109.940000 107.260000 ;
      RECT 1.000000 106.280000 109.940000 106.410000 ;
      RECT 109.210000 105.800000 109.940000 106.280000 ;
      RECT 96.560000 105.200000 107.410000 106.280000 ;
      RECT 51.560000 105.200000 94.760000 106.280000 ;
      RECT 6.560000 105.200000 49.760000 106.280000 ;
      RECT 2.530000 105.200000 4.595000 106.280000 ;
      RECT 0.000000 105.200000 0.730000 105.430000 ;
      RECT 0.000000 105.190000 108.940000 105.200000 ;
      RECT 1.000000 104.820000 108.940000 105.190000 ;
      RECT 1.000000 104.210000 109.940000 104.820000 ;
      RECT 0.000000 103.970000 109.940000 104.210000 ;
      RECT 1.000000 103.560000 109.940000 103.970000 ;
      RECT 107.410000 103.360000 109.940000 103.560000 ;
      RECT 1.000000 102.990000 2.530000 103.560000 ;
      RECT 107.410000 102.480000 108.940000 103.360000 ;
      RECT 98.560000 102.480000 105.610000 103.560000 ;
      RECT 53.560000 102.480000 96.760000 103.560000 ;
      RECT 8.560000 102.480000 51.760000 103.560000 ;
      RECT 4.330000 102.480000 6.760000 103.560000 ;
      RECT 0.000000 102.480000 2.530000 102.990000 ;
      RECT 0.000000 102.380000 108.940000 102.480000 ;
      RECT 0.000000 102.140000 109.940000 102.380000 ;
      RECT 1.000000 101.160000 109.940000 102.140000 ;
      RECT 0.000000 100.920000 109.940000 101.160000 ;
      RECT 1.000000 100.840000 108.940000 100.920000 ;
      RECT 109.210000 99.760000 109.940000 99.940000 ;
      RECT 96.560000 99.760000 107.410000 100.840000 ;
      RECT 51.560000 99.760000 94.760000 100.840000 ;
      RECT 6.560000 99.760000 49.760000 100.840000 ;
      RECT 2.530000 99.760000 4.595000 100.840000 ;
      RECT 0.000000 99.760000 0.730000 99.940000 ;
      RECT 0.000000 99.090000 109.940000 99.760000 ;
      RECT 1.000000 98.120000 108.940000 99.090000 ;
      RECT 107.410000 98.110000 108.940000 98.120000 ;
      RECT 1.000000 98.110000 2.530000 98.120000 ;
      RECT 0.000000 97.870000 2.530000 98.110000 ;
      RECT 107.410000 97.040000 109.940000 98.110000 ;
      RECT 98.560000 97.040000 105.610000 98.120000 ;
      RECT 53.560000 97.040000 96.760000 98.120000 ;
      RECT 8.560000 97.040000 51.760000 98.120000 ;
      RECT 4.330000 97.040000 6.760000 98.120000 ;
      RECT 1.000000 97.040000 2.530000 97.870000 ;
      RECT 1.000000 96.890000 109.940000 97.040000 ;
      RECT 0.000000 96.650000 109.940000 96.890000 ;
      RECT 0.000000 96.040000 108.940000 96.650000 ;
      RECT 1.000000 95.670000 108.940000 96.040000 ;
      RECT 1.000000 95.400000 109.940000 95.670000 ;
      RECT 0.000000 94.820000 0.730000 95.060000 ;
      RECT 109.210000 94.320000 109.940000 95.400000 ;
      RECT 96.560000 94.320000 107.410000 95.400000 ;
      RECT 51.560000 94.320000 94.760000 95.400000 ;
      RECT 6.560000 94.320000 49.760000 95.400000 ;
      RECT 2.530000 94.320000 4.595000 95.400000 ;
      RECT 1.000000 94.210000 109.940000 94.320000 ;
      RECT 1.000000 93.840000 108.940000 94.210000 ;
      RECT 0.000000 93.600000 108.940000 93.840000 ;
      RECT 1.000000 93.230000 108.940000 93.600000 ;
      RECT 1.000000 92.680000 109.940000 93.230000 ;
      RECT 1.000000 92.620000 2.530000 92.680000 ;
      RECT 107.410000 91.770000 109.940000 92.680000 ;
      RECT 0.000000 91.770000 2.530000 92.620000 ;
      RECT 107.410000 91.600000 108.940000 91.770000 ;
      RECT 98.560000 91.600000 105.610000 92.680000 ;
      RECT 53.560000 91.600000 96.760000 92.680000 ;
      RECT 8.560000 91.600000 51.760000 92.680000 ;
      RECT 4.330000 91.600000 6.760000 92.680000 ;
      RECT 1.000000 91.600000 2.530000 91.770000 ;
      RECT 1.000000 90.790000 108.940000 91.600000 ;
      RECT 0.000000 90.550000 109.940000 90.790000 ;
      RECT 1.000000 89.960000 109.940000 90.550000 ;
      RECT 109.210000 89.330000 109.940000 89.960000 ;
      RECT 96.560000 88.880000 107.410000 89.960000 ;
      RECT 51.560000 88.880000 94.760000 89.960000 ;
      RECT 6.560000 88.880000 49.760000 89.960000 ;
      RECT 2.530000 88.880000 4.595000 89.960000 ;
      RECT 0.000000 88.880000 0.730000 89.570000 ;
      RECT 0.000000 88.720000 108.940000 88.880000 ;
      RECT 1.000000 88.350000 108.940000 88.720000 ;
      RECT 1.000000 87.740000 109.940000 88.350000 ;
      RECT 0.000000 87.500000 109.940000 87.740000 ;
      RECT 1.000000 87.240000 109.940000 87.500000 ;
      RECT 107.410000 86.890000 109.940000 87.240000 ;
      RECT 1.000000 86.520000 2.530000 87.240000 ;
      RECT 107.410000 86.160000 108.940000 86.890000 ;
      RECT 98.560000 86.160000 105.610000 87.240000 ;
      RECT 53.560000 86.160000 96.760000 87.240000 ;
      RECT 8.560000 86.160000 51.760000 87.240000 ;
      RECT 4.330000 86.160000 6.760000 87.240000 ;
      RECT 0.000000 86.160000 2.530000 86.520000 ;
      RECT 0.000000 85.910000 108.940000 86.160000 ;
      RECT 0.000000 85.670000 109.940000 85.910000 ;
      RECT 1.000000 84.690000 109.940000 85.670000 ;
      RECT 0.000000 84.520000 109.940000 84.690000 ;
      RECT 109.210000 84.450000 109.940000 84.520000 ;
      RECT 0.000000 84.450000 0.730000 84.520000 ;
      RECT 109.210000 83.440000 109.940000 83.470000 ;
      RECT 96.560000 83.440000 107.410000 84.520000 ;
      RECT 51.560000 83.440000 94.760000 84.520000 ;
      RECT 6.560000 83.440000 49.760000 84.520000 ;
      RECT 2.530000 83.440000 4.595000 84.520000 ;
      RECT 0.000000 83.440000 0.730000 83.470000 ;
      RECT 0.000000 82.620000 109.940000 83.440000 ;
      RECT 1.000000 82.010000 109.940000 82.620000 ;
      RECT 1.000000 81.800000 108.940000 82.010000 ;
      RECT 1.000000 81.640000 2.530000 81.800000 ;
      RECT 0.000000 81.400000 2.530000 81.640000 ;
      RECT 107.410000 81.030000 108.940000 81.800000 ;
      RECT 107.410000 80.720000 109.940000 81.030000 ;
      RECT 98.560000 80.720000 105.610000 81.800000 ;
      RECT 53.560000 80.720000 96.760000 81.800000 ;
      RECT 8.560000 80.720000 51.760000 81.800000 ;
      RECT 4.330000 80.720000 6.760000 81.800000 ;
      RECT 1.000000 80.720000 2.530000 81.400000 ;
      RECT 1.000000 80.420000 109.940000 80.720000 ;
      RECT 0.000000 80.180000 109.940000 80.420000 ;
      RECT 1.000000 79.570000 109.940000 80.180000 ;
      RECT 1.000000 79.200000 108.940000 79.570000 ;
      RECT 0.000000 79.080000 108.940000 79.200000 ;
      RECT 0.000000 78.350000 0.730000 79.080000 ;
      RECT 109.210000 78.000000 109.940000 78.590000 ;
      RECT 96.560000 78.000000 107.410000 79.080000 ;
      RECT 51.560000 78.000000 94.760000 79.080000 ;
      RECT 6.560000 78.000000 49.760000 79.080000 ;
      RECT 2.530000 78.000000 4.595000 79.080000 ;
      RECT 1.000000 77.370000 109.940000 78.000000 ;
      RECT 0.000000 77.130000 109.940000 77.370000 ;
      RECT 1.000000 76.360000 108.940000 77.130000 ;
      RECT 107.410000 76.150000 108.940000 76.360000 ;
      RECT 1.000000 76.150000 2.530000 76.360000 ;
      RECT 0.000000 75.300000 2.530000 76.150000 ;
      RECT 107.410000 75.280000 109.940000 76.150000 ;
      RECT 98.560000 75.280000 105.610000 76.360000 ;
      RECT 53.560000 75.280000 96.760000 76.360000 ;
      RECT 8.560000 75.280000 51.760000 76.360000 ;
      RECT 4.330000 75.280000 6.760000 76.360000 ;
      RECT 1.000000 75.280000 2.530000 75.300000 ;
      RECT 1.000000 74.690000 109.940000 75.280000 ;
      RECT 1.000000 74.320000 108.940000 74.690000 ;
      RECT 0.000000 74.080000 108.940000 74.320000 ;
      RECT 1.000000 73.710000 108.940000 74.080000 ;
      RECT 1.000000 73.640000 109.940000 73.710000 ;
      RECT 109.210000 72.560000 109.940000 73.640000 ;
      RECT 96.560000 72.560000 107.410000 73.640000 ;
      RECT 51.560000 72.560000 94.760000 73.640000 ;
      RECT 6.560000 72.560000 49.760000 73.640000 ;
      RECT 2.530000 72.560000 4.595000 73.640000 ;
      RECT 0.000000 72.560000 0.730000 73.100000 ;
      RECT 0.000000 72.250000 109.940000 72.560000 ;
      RECT 1.000000 71.270000 108.940000 72.250000 ;
      RECT 0.000000 71.030000 109.940000 71.270000 ;
      RECT 1.000000 70.920000 109.940000 71.030000 ;
      RECT 1.000000 70.050000 2.530000 70.920000 ;
      RECT 107.410000 69.840000 109.940000 70.920000 ;
      RECT 98.560000 69.840000 105.610000 70.920000 ;
      RECT 53.560000 69.840000 96.760000 70.920000 ;
      RECT 8.560000 69.840000 51.760000 70.920000 ;
      RECT 4.330000 69.840000 6.760000 70.920000 ;
      RECT 0.000000 69.840000 2.530000 70.050000 ;
      RECT 0.000000 69.810000 109.940000 69.840000 ;
      RECT 0.000000 69.200000 108.940000 69.810000 ;
      RECT 1.000000 68.830000 108.940000 69.200000 ;
      RECT 1.000000 68.220000 109.940000 68.830000 ;
      RECT 0.000000 68.200000 109.940000 68.220000 ;
      RECT 109.210000 67.980000 109.940000 68.200000 ;
      RECT 0.000000 67.980000 0.730000 68.200000 ;
      RECT 96.560000 67.120000 107.410000 68.200000 ;
      RECT 51.560000 67.120000 94.760000 68.200000 ;
      RECT 6.560000 67.120000 49.760000 68.200000 ;
      RECT 2.530000 67.120000 4.595000 68.200000 ;
      RECT 1.000000 67.000000 108.940000 67.120000 ;
      RECT 0.000000 66.760000 109.940000 67.000000 ;
      RECT 1.000000 65.780000 109.940000 66.760000 ;
      RECT 0.000000 65.540000 109.940000 65.780000 ;
      RECT 0.000000 65.480000 108.940000 65.540000 ;
      RECT 0.000000 64.930000 2.530000 65.480000 ;
      RECT 107.410000 64.560000 108.940000 65.480000 ;
      RECT 107.410000 64.400000 109.940000 64.560000 ;
      RECT 98.560000 64.400000 105.610000 65.480000 ;
      RECT 53.560000 64.400000 96.760000 65.480000 ;
      RECT 8.560000 64.400000 51.760000 65.480000 ;
      RECT 4.330000 64.400000 6.760000 65.480000 ;
      RECT 1.000000 64.400000 2.530000 64.930000 ;
      RECT 1.000000 63.950000 109.940000 64.400000 ;
      RECT 0.000000 63.710000 109.940000 63.950000 ;
      RECT 1.000000 63.100000 109.940000 63.710000 ;
      RECT 1.000000 62.760000 108.940000 63.100000 ;
      RECT 0.000000 61.880000 0.730000 62.730000 ;
      RECT 109.210000 61.680000 109.940000 62.120000 ;
      RECT 96.560000 61.680000 107.410000 62.760000 ;
      RECT 51.560000 61.680000 94.760000 62.760000 ;
      RECT 6.560000 61.680000 49.760000 62.760000 ;
      RECT 2.530000 61.680000 4.595000 62.760000 ;
      RECT 1.000000 60.900000 109.940000 61.680000 ;
      RECT 0.000000 60.660000 109.940000 60.900000 ;
      RECT 1.000000 60.040000 108.940000 60.660000 ;
      RECT 107.410000 59.680000 108.940000 60.040000 ;
      RECT 1.000000 59.680000 2.530000 60.040000 ;
      RECT 107.410000 58.960000 109.940000 59.680000 ;
      RECT 98.560000 58.960000 105.610000 60.040000 ;
      RECT 53.560000 58.960000 96.760000 60.040000 ;
      RECT 8.560000 58.960000 51.760000 60.040000 ;
      RECT 4.330000 58.960000 6.760000 60.040000 ;
      RECT 0.000000 58.960000 2.530000 59.680000 ;
      RECT 0.000000 58.830000 109.940000 58.960000 ;
      RECT 1.000000 58.220000 109.940000 58.830000 ;
      RECT 1.000000 57.850000 108.940000 58.220000 ;
      RECT 0.000000 57.610000 108.940000 57.850000 ;
      RECT 1.000000 57.320000 108.940000 57.610000 ;
      RECT 109.210000 56.240000 109.940000 57.240000 ;
      RECT 96.560000 56.240000 107.410000 57.320000 ;
      RECT 51.560000 56.240000 94.760000 57.320000 ;
      RECT 6.560000 56.240000 49.760000 57.320000 ;
      RECT 2.530000 56.240000 4.595000 57.320000 ;
      RECT 0.000000 56.240000 0.730000 56.630000 ;
      RECT 0.000000 55.780000 109.940000 56.240000 ;
      RECT 1.000000 54.800000 108.940000 55.780000 ;
      RECT 0.000000 54.600000 109.940000 54.800000 ;
      RECT 0.000000 54.560000 2.530000 54.600000 ;
      RECT 1.000000 53.580000 2.530000 54.560000 ;
      RECT 107.410000 53.520000 109.940000 54.600000 ;
      RECT 98.560000 53.520000 105.610000 54.600000 ;
      RECT 53.560000 53.520000 96.760000 54.600000 ;
      RECT 8.560000 53.520000 51.760000 54.600000 ;
      RECT 4.330000 53.520000 6.760000 54.600000 ;
      RECT 0.000000 53.520000 2.530000 53.580000 ;
      RECT 0.000000 53.340000 109.940000 53.520000 ;
      RECT 1.000000 52.360000 108.940000 53.340000 ;
      RECT 0.000000 51.880000 109.940000 52.360000 ;
      RECT 0.000000 51.510000 0.730000 51.880000 ;
      RECT 109.210000 50.900000 109.940000 51.880000 ;
      RECT 96.560000 50.800000 107.410000 51.880000 ;
      RECT 51.560000 50.800000 94.760000 51.880000 ;
      RECT 6.560000 50.800000 49.760000 51.880000 ;
      RECT 2.530000 50.800000 4.595000 51.880000 ;
      RECT 1.000000 50.530000 108.940000 50.800000 ;
      RECT 0.000000 50.290000 108.940000 50.530000 ;
      RECT 1.000000 49.920000 108.940000 50.290000 ;
      RECT 1.000000 49.310000 109.940000 49.920000 ;
      RECT 0.000000 49.160000 109.940000 49.310000 ;
      RECT 107.410000 48.460000 109.940000 49.160000 ;
      RECT 0.000000 48.460000 2.530000 49.160000 ;
      RECT 107.410000 48.080000 108.940000 48.460000 ;
      RECT 98.560000 48.080000 105.610000 49.160000 ;
      RECT 53.560000 48.080000 96.760000 49.160000 ;
      RECT 8.560000 48.080000 51.760000 49.160000 ;
      RECT 4.330000 48.080000 6.760000 49.160000 ;
      RECT 1.000000 48.080000 2.530000 48.460000 ;
      RECT 1.000000 47.480000 108.940000 48.080000 ;
      RECT 0.000000 47.240000 109.940000 47.480000 ;
      RECT 1.000000 46.440000 109.940000 47.240000 ;
      RECT 109.210000 46.020000 109.940000 46.440000 ;
      RECT 0.000000 45.410000 0.730000 46.260000 ;
      RECT 96.560000 45.360000 107.410000 46.440000 ;
      RECT 51.560000 45.360000 94.760000 46.440000 ;
      RECT 6.560000 45.360000 49.760000 46.440000 ;
      RECT 2.530000 45.360000 4.595000 46.440000 ;
      RECT 1.000000 45.040000 108.940000 45.360000 ;
      RECT 1.000000 44.430000 109.940000 45.040000 ;
      RECT 0.000000 44.190000 109.940000 44.430000 ;
      RECT 1.000000 43.720000 109.940000 44.190000 ;
      RECT 107.410000 43.580000 109.940000 43.720000 ;
      RECT 1.000000 43.210000 2.530000 43.720000 ;
      RECT 0.000000 42.970000 2.530000 43.210000 ;
      RECT 107.410000 42.640000 108.940000 43.580000 ;
      RECT 98.560000 42.640000 105.610000 43.720000 ;
      RECT 53.560000 42.640000 96.760000 43.720000 ;
      RECT 8.560000 42.640000 51.760000 43.720000 ;
      RECT 4.330000 42.640000 6.760000 43.720000 ;
      RECT 1.000000 42.640000 2.530000 42.970000 ;
      RECT 1.000000 42.600000 108.940000 42.640000 ;
      RECT 1.000000 41.990000 109.940000 42.600000 ;
      RECT 0.000000 41.140000 109.940000 41.990000 ;
      RECT 1.000000 41.000000 108.940000 41.140000 ;
      RECT 109.210000 39.920000 109.940000 40.160000 ;
      RECT 96.560000 39.920000 107.410000 41.000000 ;
      RECT 51.560000 39.920000 94.760000 41.000000 ;
      RECT 6.560000 39.920000 49.760000 41.000000 ;
      RECT 2.530000 39.920000 4.595000 41.000000 ;
      RECT 0.000000 39.920000 0.730000 40.160000 ;
      RECT 1.000000 38.940000 109.940000 39.920000 ;
      RECT 0.000000 38.700000 109.940000 38.940000 ;
      RECT 0.000000 38.280000 108.940000 38.700000 ;
      RECT 0.000000 38.090000 2.530000 38.280000 ;
      RECT 107.410000 37.720000 108.940000 38.280000 ;
      RECT 107.410000 37.200000 109.940000 37.720000 ;
      RECT 98.560000 37.200000 105.610000 38.280000 ;
      RECT 53.560000 37.200000 96.760000 38.280000 ;
      RECT 8.560000 37.200000 51.760000 38.280000 ;
      RECT 4.330000 37.200000 6.760000 38.280000 ;
      RECT 1.000000 37.200000 2.530000 38.090000 ;
      RECT 1.000000 37.110000 109.940000 37.200000 ;
      RECT 0.000000 36.870000 109.940000 37.110000 ;
      RECT 1.000000 35.890000 108.940000 36.870000 ;
      RECT 0.000000 35.560000 109.940000 35.890000 ;
      RECT 0.000000 35.040000 0.730000 35.560000 ;
      RECT 109.210000 34.480000 109.940000 35.560000 ;
      RECT 96.560000 34.480000 107.410000 35.560000 ;
      RECT 51.560000 34.480000 94.760000 35.560000 ;
      RECT 6.560000 34.480000 49.760000 35.560000 ;
      RECT 2.530000 34.480000 4.595000 35.560000 ;
      RECT 1.000000 34.430000 109.940000 34.480000 ;
      RECT 1.000000 34.060000 108.940000 34.430000 ;
      RECT 0.000000 33.820000 108.940000 34.060000 ;
      RECT 1.000000 33.450000 108.940000 33.820000 ;
      RECT 1.000000 32.840000 109.940000 33.450000 ;
      RECT 107.410000 31.990000 109.940000 32.840000 ;
      RECT 0.000000 31.990000 2.530000 32.840000 ;
      RECT 107.410000 31.760000 108.940000 31.990000 ;
      RECT 98.560000 31.760000 105.610000 32.840000 ;
      RECT 53.560000 31.760000 96.760000 32.840000 ;
      RECT 8.560000 31.760000 51.760000 32.840000 ;
      RECT 4.330000 31.760000 6.760000 32.840000 ;
      RECT 1.000000 31.760000 2.530000 31.990000 ;
      RECT 1.000000 31.010000 108.940000 31.760000 ;
      RECT 0.000000 30.770000 109.940000 31.010000 ;
      RECT 1.000000 30.120000 109.940000 30.770000 ;
      RECT 109.210000 29.550000 109.940000 30.120000 ;
      RECT 0.000000 29.550000 0.730000 29.790000 ;
      RECT 96.560000 29.040000 107.410000 30.120000 ;
      RECT 51.560000 29.040000 94.760000 30.120000 ;
      RECT 6.560000 29.040000 49.760000 30.120000 ;
      RECT 2.530000 29.040000 4.595000 30.120000 ;
      RECT 1.000000 28.570000 108.940000 29.040000 ;
      RECT 0.000000 27.720000 109.940000 28.570000 ;
      RECT 1.000000 27.400000 109.940000 27.720000 ;
      RECT 107.410000 27.110000 109.940000 27.400000 ;
      RECT 1.000000 26.740000 2.530000 27.400000 ;
      RECT 0.000000 26.500000 2.530000 26.740000 ;
      RECT 107.410000 26.320000 108.940000 27.110000 ;
      RECT 98.560000 26.320000 105.610000 27.400000 ;
      RECT 53.560000 26.320000 96.760000 27.400000 ;
      RECT 8.560000 26.320000 51.760000 27.400000 ;
      RECT 4.330000 26.320000 6.760000 27.400000 ;
      RECT 1.000000 26.320000 2.530000 26.500000 ;
      RECT 1.000000 26.130000 108.940000 26.320000 ;
      RECT 1.000000 25.520000 109.940000 26.130000 ;
      RECT 0.000000 24.680000 109.940000 25.520000 ;
      RECT 109.210000 24.670000 109.940000 24.680000 ;
      RECT 0.000000 24.670000 0.730000 24.680000 ;
      RECT 109.210000 23.600000 109.940000 23.690000 ;
      RECT 96.560000 23.600000 107.410000 24.680000 ;
      RECT 51.560000 23.600000 94.760000 24.680000 ;
      RECT 6.560000 23.600000 49.760000 24.680000 ;
      RECT 2.530000 23.600000 4.595000 24.680000 ;
      RECT 0.000000 23.600000 0.730000 23.690000 ;
      RECT 0.000000 23.450000 109.940000 23.600000 ;
      RECT 1.000000 22.470000 109.940000 23.450000 ;
      RECT 0.000000 22.230000 109.940000 22.470000 ;
      RECT 0.000000 21.960000 108.940000 22.230000 ;
      RECT 0.000000 21.620000 2.530000 21.960000 ;
      RECT 107.410000 21.250000 108.940000 21.960000 ;
      RECT 107.410000 20.880000 109.940000 21.250000 ;
      RECT 98.560000 20.880000 105.610000 21.960000 ;
      RECT 53.560000 20.880000 96.760000 21.960000 ;
      RECT 8.560000 20.880000 51.760000 21.960000 ;
      RECT 4.330000 20.880000 6.760000 21.960000 ;
      RECT 1.000000 20.880000 2.530000 21.620000 ;
      RECT 1.000000 20.640000 109.940000 20.880000 ;
      RECT 0.000000 20.400000 109.940000 20.640000 ;
      RECT 1.000000 19.790000 109.940000 20.400000 ;
      RECT 1.000000 19.420000 108.940000 19.790000 ;
      RECT 0.000000 19.240000 108.940000 19.420000 ;
      RECT 0.000000 18.570000 0.730000 19.240000 ;
      RECT 109.210000 18.160000 109.940000 18.810000 ;
      RECT 96.560000 18.160000 107.410000 19.240000 ;
      RECT 51.560000 18.160000 94.760000 19.240000 ;
      RECT 6.560000 18.160000 49.760000 19.240000 ;
      RECT 2.530000 18.160000 4.595000 19.240000 ;
      RECT 1.000000 17.590000 109.940000 18.160000 ;
      RECT 0.000000 17.350000 109.940000 17.590000 ;
      RECT 1.000000 16.520000 108.940000 17.350000 ;
      RECT 107.410000 16.370000 108.940000 16.520000 ;
      RECT 1.000000 16.370000 2.530000 16.520000 ;
      RECT 0.000000 16.130000 2.530000 16.370000 ;
      RECT 107.410000 15.440000 109.940000 16.370000 ;
      RECT 98.560000 15.440000 105.610000 16.520000 ;
      RECT 53.560000 15.440000 96.760000 16.520000 ;
      RECT 8.560000 15.440000 51.760000 16.520000 ;
      RECT 4.330000 15.440000 6.760000 16.520000 ;
      RECT 1.000000 15.440000 2.530000 16.130000 ;
      RECT 1.000000 15.150000 109.940000 15.440000 ;
      RECT 0.000000 14.910000 109.940000 15.150000 ;
      RECT 0.000000 14.300000 108.940000 14.910000 ;
      RECT 1.000000 13.930000 108.940000 14.300000 ;
      RECT 1.000000 13.800000 109.940000 13.930000 ;
      RECT 0.000000 13.080000 0.730000 13.320000 ;
      RECT 109.210000 12.720000 109.940000 13.800000 ;
      RECT 96.560000 12.720000 107.410000 13.800000 ;
      RECT 51.560000 12.720000 94.760000 13.800000 ;
      RECT 6.560000 12.720000 49.760000 13.800000 ;
      RECT 2.530000 12.720000 4.595000 13.800000 ;
      RECT 1.000000 12.470000 109.940000 12.720000 ;
      RECT 1.000000 12.100000 108.940000 12.470000 ;
      RECT 0.000000 11.490000 108.940000 12.100000 ;
      RECT 0.000000 11.250000 109.940000 11.490000 ;
      RECT 1.000000 11.080000 109.940000 11.250000 ;
      RECT 1.000000 10.270000 2.530000 11.080000 ;
      RECT 107.410000 10.030000 109.940000 11.080000 ;
      RECT 0.000000 10.030000 2.530000 10.270000 ;
      RECT 107.410000 10.000000 108.940000 10.030000 ;
      RECT 98.560000 10.000000 105.610000 11.080000 ;
      RECT 53.560000 10.000000 96.760000 11.080000 ;
      RECT 8.560000 10.000000 51.760000 11.080000 ;
      RECT 4.330000 10.000000 6.760000 11.080000 ;
      RECT 1.000000 10.000000 2.530000 10.030000 ;
      RECT 1.000000 9.050000 108.940000 10.000000 ;
      RECT 0.000000 8.360000 109.940000 9.050000 ;
      RECT 0.000000 8.200000 0.730000 8.360000 ;
      RECT 109.210000 7.590000 109.940000 8.360000 ;
      RECT 96.560000 7.280000 107.410000 8.360000 ;
      RECT 51.560000 7.280000 94.760000 8.360000 ;
      RECT 6.560000 7.280000 49.760000 8.360000 ;
      RECT 2.530000 7.280000 4.595000 8.360000 ;
      RECT 1.000000 7.220000 108.940000 7.280000 ;
      RECT 0.000000 6.980000 108.940000 7.220000 ;
      RECT 1.000000 6.610000 108.940000 6.980000 ;
      RECT 1.000000 6.000000 109.940000 6.610000 ;
      RECT 0.000000 5.760000 109.940000 6.000000 ;
      RECT 1.000000 5.640000 108.940000 5.760000 ;
      RECT 107.410000 4.780000 108.940000 5.640000 ;
      RECT 1.000000 4.780000 2.530000 5.640000 ;
      RECT 107.410000 4.560000 109.940000 4.780000 ;
      RECT 98.560000 4.560000 105.610000 5.640000 ;
      RECT 53.560000 4.560000 96.760000 5.640000 ;
      RECT 8.560000 4.560000 51.760000 5.640000 ;
      RECT 4.330000 4.560000 6.760000 5.640000 ;
      RECT 0.000000 4.560000 2.530000 4.780000 ;
      RECT 0.000000 4.350000 109.940000 4.560000 ;
      RECT 0.000000 0.000000 109.940000 0.750000 ;
    LAYER met4 ;
      RECT 4.330000 198.320000 105.610000 200.260000 ;
      RECT 96.560000 196.520000 105.610000 198.320000 ;
      RECT 51.560000 196.520000 94.760000 198.320000 ;
      RECT 6.560000 196.520000 49.760000 198.320000 ;
      RECT 4.330000 193.320000 4.760000 198.320000 ;
      RECT 4.330000 192.240000 4.595000 193.320000 ;
      RECT 4.330000 187.880000 4.760000 192.240000 ;
      RECT 4.330000 186.800000 4.595000 187.880000 ;
      RECT 4.330000 182.440000 4.760000 186.800000 ;
      RECT 4.330000 181.360000 4.595000 182.440000 ;
      RECT 4.330000 177.000000 4.760000 181.360000 ;
      RECT 4.330000 175.920000 4.595000 177.000000 ;
      RECT 4.330000 171.560000 4.760000 175.920000 ;
      RECT 4.330000 170.480000 4.595000 171.560000 ;
      RECT 4.330000 166.120000 4.760000 170.480000 ;
      RECT 4.330000 165.040000 4.595000 166.120000 ;
      RECT 4.330000 160.680000 4.760000 165.040000 ;
      RECT 4.330000 159.600000 4.595000 160.680000 ;
      RECT 4.330000 155.240000 4.760000 159.600000 ;
      RECT 4.330000 154.160000 4.595000 155.240000 ;
      RECT 4.330000 149.800000 4.760000 154.160000 ;
      RECT 4.330000 148.720000 4.595000 149.800000 ;
      RECT 4.330000 144.360000 4.760000 148.720000 ;
      RECT 4.330000 143.280000 4.595000 144.360000 ;
      RECT 4.330000 138.920000 4.760000 143.280000 ;
      RECT 4.330000 137.840000 4.595000 138.920000 ;
      RECT 4.330000 133.480000 4.760000 137.840000 ;
      RECT 4.330000 132.400000 4.595000 133.480000 ;
      RECT 4.330000 128.040000 4.760000 132.400000 ;
      RECT 4.330000 126.960000 4.595000 128.040000 ;
      RECT 4.330000 122.600000 4.760000 126.960000 ;
      RECT 4.330000 121.520000 4.595000 122.600000 ;
      RECT 4.330000 117.160000 4.760000 121.520000 ;
      RECT 4.330000 116.080000 4.595000 117.160000 ;
      RECT 4.330000 111.720000 4.760000 116.080000 ;
      RECT 4.330000 110.640000 4.595000 111.720000 ;
      RECT 4.330000 106.280000 4.760000 110.640000 ;
      RECT 4.330000 105.200000 4.595000 106.280000 ;
      RECT 4.330000 100.840000 4.760000 105.200000 ;
      RECT 4.330000 99.760000 4.595000 100.840000 ;
      RECT 4.330000 95.400000 4.760000 99.760000 ;
      RECT 4.330000 94.320000 4.595000 95.400000 ;
      RECT 4.330000 89.960000 4.760000 94.320000 ;
      RECT 4.330000 88.880000 4.595000 89.960000 ;
      RECT 4.330000 84.520000 4.760000 88.880000 ;
      RECT 4.330000 83.440000 4.595000 84.520000 ;
      RECT 4.330000 79.080000 4.760000 83.440000 ;
      RECT 4.330000 78.000000 4.595000 79.080000 ;
      RECT 4.330000 73.640000 4.760000 78.000000 ;
      RECT 4.330000 72.560000 4.595000 73.640000 ;
      RECT 4.330000 68.200000 4.760000 72.560000 ;
      RECT 4.330000 67.120000 4.595000 68.200000 ;
      RECT 4.330000 62.760000 4.760000 67.120000 ;
      RECT 4.330000 61.680000 4.595000 62.760000 ;
      RECT 4.330000 57.320000 4.760000 61.680000 ;
      RECT 4.330000 56.240000 4.595000 57.320000 ;
      RECT 4.330000 51.880000 4.760000 56.240000 ;
      RECT 4.330000 50.800000 4.595000 51.880000 ;
      RECT 4.330000 46.440000 4.760000 50.800000 ;
      RECT 4.330000 45.360000 4.595000 46.440000 ;
      RECT 4.330000 41.000000 4.760000 45.360000 ;
      RECT 4.330000 39.920000 4.595000 41.000000 ;
      RECT 4.330000 35.560000 4.760000 39.920000 ;
      RECT 4.330000 34.480000 4.595000 35.560000 ;
      RECT 4.330000 30.120000 4.760000 34.480000 ;
      RECT 4.330000 29.040000 4.595000 30.120000 ;
      RECT 4.330000 24.680000 4.760000 29.040000 ;
      RECT 4.330000 23.600000 4.595000 24.680000 ;
      RECT 4.330000 19.240000 4.760000 23.600000 ;
      RECT 4.330000 18.160000 4.595000 19.240000 ;
      RECT 4.330000 13.800000 4.760000 18.160000 ;
      RECT 4.330000 12.720000 4.595000 13.800000 ;
      RECT 4.330000 8.360000 4.760000 12.720000 ;
      RECT 4.330000 7.280000 4.595000 8.360000 ;
      RECT 98.560000 2.550000 105.610000 196.520000 ;
      RECT 96.560000 2.550000 96.760000 196.520000 ;
      RECT 53.560000 2.550000 94.760000 196.520000 ;
      RECT 51.560000 2.550000 51.760000 196.520000 ;
      RECT 8.560000 2.550000 49.760000 196.520000 ;
      RECT 6.560000 2.550000 6.760000 196.520000 ;
      RECT 96.560000 0.750000 105.610000 2.550000 ;
      RECT 51.560000 0.750000 94.760000 2.550000 ;
      RECT 6.560000 0.750000 49.760000 2.550000 ;
      RECT 4.330000 0.750000 4.760000 7.280000 ;
      RECT 109.210000 0.000000 109.940000 200.260000 ;
      RECT 4.330000 0.000000 105.610000 0.750000 ;
      RECT 0.000000 0.000000 0.730000 200.260000 ;
  END
END RAM_IO

END LIBRARY
